-- Input HEX file name : test_fix_fft.ihex
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity programToLoad is port (
address_in : in  std_logic_vector (15 downto 0);
data_out   : out std_logic_vector (15 downto 0));
end programToLoad;

architecture rtl of programToLoad is
begin
data_out <=
		x"940C" when address_in = 16#0000# else
		x"0430" when address_in = 16#0001# else
		x"940C" when address_in = 16#0002# else
		x"0450" when address_in = 16#0003# else
		x"940C" when address_in = 16#0004# else
		x"0450" when address_in = 16#0005# else
		x"940C" when address_in = 16#0006# else
		x"0450" when address_in = 16#0007# else
		x"940C" when address_in = 16#0008# else
		x"0450" when address_in = 16#0009# else
		x"940C" when address_in = 16#000A# else
		x"0450" when address_in = 16#000B# else
		x"940C" when address_in = 16#000C# else
		x"0450" when address_in = 16#000D# else
		x"940C" when address_in = 16#000E# else
		x"0450" when address_in = 16#000F# else
		x"940C" when address_in = 16#0010# else
		x"0450" when address_in = 16#0011# else
		x"940C" when address_in = 16#0012# else
		x"0450" when address_in = 16#0013# else
		x"940C" when address_in = 16#0014# else
		x"0450" when address_in = 16#0015# else
		x"940C" when address_in = 16#0016# else
		x"0450" when address_in = 16#0017# else
		x"940C" when address_in = 16#0018# else
		x"0450" when address_in = 16#0019# else
		x"940C" when address_in = 16#001A# else
		x"0450" when address_in = 16#001B# else
		x"940C" when address_in = 16#001C# else
		x"0450" when address_in = 16#001D# else
		x"940C" when address_in = 16#001E# else
		x"0450" when address_in = 16#001F# else
		x"940C" when address_in = 16#0020# else
		x"0450" when address_in = 16#0021# else
		x"940C" when address_in = 16#0022# else
		x"0450" when address_in = 16#0023# else
		x"940C" when address_in = 16#0024# else
		x"0450" when address_in = 16#0025# else
		x"940C" when address_in = 16#0026# else
		x"0450" when address_in = 16#0027# else
		x"940C" when address_in = 16#0028# else
		x"0450" when address_in = 16#0029# else
		x"940C" when address_in = 16#002A# else
		x"0450" when address_in = 16#002B# else
		x"940C" when address_in = 16#002C# else
		x"0450" when address_in = 16#002D# else
		x"940C" when address_in = 16#002E# else
		x"0450" when address_in = 16#002F# else
		x"3000" when address_in = 16#0030# else
		x"2FA3" when address_in = 16#0031# else
		x"2E8F" when address_in = 16#0032# else
		x"2CC8" when address_in = 16#0033# else
		x"2A55" when address_in = 16#0034# else
		x"273E" when address_in = 16#0035# else
		x"2390" when address_in = 16#0036# else
		x"1F5A" when address_in = 16#0037# else
		x"1AAA" when address_in = 16#0038# else
		x"1594" when address_in = 16#0039# else
		x"102B" when address_in = 16#003A# else
		x"0A84" when address_in = 16#003B# else
		x"04B4" when address_in = 16#003C# else
		x"FED3" when address_in = 16#003D# else
		x"F8F5" when address_in = 16#003E# else
		x"F333" when address_in = 16#003F# else
		x"EDA2" when address_in = 16#0040# else
		x"E858" when address_in = 16#0041# else
		x"E369" when address_in = 16#0042# else
		x"DEE7" when address_in = 16#0043# else
		x"DAE6" when address_in = 16#0044# else
		x"D773" when address_in = 16#0045# else
		x"D49C" when address_in = 16#0046# else
		x"D26D" when address_in = 16#0047# else
		x"D0ED" when address_in = 16#0048# else
		x"D022" when address_in = 16#0049# else
		x"D00F" when address_in = 16#004A# else
		x"D0B5" when address_in = 16#004B# else
		x"D212" when address_in = 16#004C# else
		x"D41F" when address_in = 16#004D# else
		x"D6D5" when address_in = 16#004E# else
		x"DA29" when address_in = 16#004F# else
		x"DE10" when address_in = 16#0050# else
		x"E279" when address_in = 16#0051# else
		x"E753" when address_in = 16#0052# else
		x"EC8D" when address_in = 16#0053# else
		x"F211" when address_in = 16#0054# else
		x"F7CC" when address_in = 16#0055# else
		x"FDA6" when address_in = 16#0056# else
		x"0387" when address_in = 16#0057# else
		x"095D" when address_in = 16#0058# else
		x"0F0E" when address_in = 16#0059# else
		x"1485" when address_in = 16#005A# else
		x"19AE" when address_in = 16#005B# else
		x"1E73" when address_in = 16#005C# else
		x"22C3" when address_in = 16#005D# else
		x"268D" when address_in = 16#005E# else
		x"29C3" when address_in = 16#005F# else
		x"2C58" when address_in = 16#0060# else
		x"2E42" when address_in = 16#0061# else
		x"2F7B" when address_in = 16#0062# else
		x"2FFC" when address_in = 16#0063# else
		x"2FC4" when address_in = 16#0064# else
		x"2ED5" when address_in = 16#0065# else
		x"2D31" when address_in = 16#0066# else
		x"2ADF" when address_in = 16#0067# else
		x"27E9" when address_in = 16#0068# else
		x"2458" when address_in = 16#0069# else
		x"203C" when address_in = 16#006A# else
		x"1BA3" when address_in = 16#006B# else
		x"16A0" when address_in = 16#006C# else
		x"1146" when address_in = 16#006D# else
		x"0BA9" when address_in = 16#006E# else
		x"05E0" when address_in = 16#006F# else
		x"0000" when address_in = 16#0070# else
		x"FA20" when address_in = 16#0071# else
		x"F457" when address_in = 16#0072# else
		x"EEBA" when address_in = 16#0073# else
		x"E960" when address_in = 16#0074# else
		x"E45D" when address_in = 16#0075# else
		x"DFC4" when address_in = 16#0076# else
		x"DBA8" when address_in = 16#0077# else
		x"D817" when address_in = 16#0078# else
		x"D521" when address_in = 16#0079# else
		x"D2CF" when address_in = 16#007A# else
		x"D12B" when address_in = 16#007B# else
		x"D03C" when address_in = 16#007C# else
		x"D004" when address_in = 16#007D# else
		x"D085" when address_in = 16#007E# else
		x"D1BE" when address_in = 16#007F# else
		x"D3A8" when address_in = 16#0080# else
		x"D63D" when address_in = 16#0081# else
		x"D973" when address_in = 16#0082# else
		x"DD3D" when address_in = 16#0083# else
		x"E18D" when address_in = 16#0084# else
		x"E652" when address_in = 16#0085# else
		x"EB7B" when address_in = 16#0086# else
		x"F0F2" when address_in = 16#0087# else
		x"F6A3" when address_in = 16#0088# else
		x"FC79" when address_in = 16#0089# else
		x"025A" when address_in = 16#008A# else
		x"0834" when address_in = 16#008B# else
		x"0DEF" when address_in = 16#008C# else
		x"1373" when address_in = 16#008D# else
		x"18AD" when address_in = 16#008E# else
		x"1D87" when address_in = 16#008F# else
		x"21F0" when address_in = 16#0090# else
		x"25D7" when address_in = 16#0091# else
		x"292B" when address_in = 16#0092# else
		x"2BE1" when address_in = 16#0093# else
		x"2DEE" when address_in = 16#0094# else
		x"2F4B" when address_in = 16#0095# else
		x"2FF1" when address_in = 16#0096# else
		x"2FDE" when address_in = 16#0097# else
		x"2F13" when address_in = 16#0098# else
		x"2D93" when address_in = 16#0099# else
		x"2B64" when address_in = 16#009A# else
		x"288D" when address_in = 16#009B# else
		x"251A" when address_in = 16#009C# else
		x"2119" when address_in = 16#009D# else
		x"1C97" when address_in = 16#009E# else
		x"17A8" when address_in = 16#009F# else
		x"125E" when address_in = 16#00A0# else
		x"0CCD" when address_in = 16#00A1# else
		x"070B" when address_in = 16#00A2# else
		x"012D" when address_in = 16#00A3# else
		x"FB4C" when address_in = 16#00A4# else
		x"F57C" when address_in = 16#00A5# else
		x"EFD5" when address_in = 16#00A6# else
		x"EA6C" when address_in = 16#00A7# else
		x"E556" when address_in = 16#00A8# else
		x"E0A6" when address_in = 16#00A9# else
		x"DC70" when address_in = 16#00AA# else
		x"D8C2" when address_in = 16#00AB# else
		x"D5AB" when address_in = 16#00AC# else
		x"D338" when address_in = 16#00AD# else
		x"D171" when address_in = 16#00AE# else
		x"D05D" when address_in = 16#00AF# else
		x"D000" when address_in = 16#00B0# else
		x"D05D" when address_in = 16#00B1# else
		x"D171" when address_in = 16#00B2# else
		x"D338" when address_in = 16#00B3# else
		x"D5AB" when address_in = 16#00B4# else
		x"D8C2" when address_in = 16#00B5# else
		x"DC70" when address_in = 16#00B6# else
		x"E0A6" when address_in = 16#00B7# else
		x"E556" when address_in = 16#00B8# else
		x"EA6C" when address_in = 16#00B9# else
		x"EFD5" when address_in = 16#00BA# else
		x"F57C" when address_in = 16#00BB# else
		x"FB4C" when address_in = 16#00BC# else
		x"012D" when address_in = 16#00BD# else
		x"070B" when address_in = 16#00BE# else
		x"0CCD" when address_in = 16#00BF# else
		x"125E" when address_in = 16#00C0# else
		x"17A8" when address_in = 16#00C1# else
		x"1C97" when address_in = 16#00C2# else
		x"2119" when address_in = 16#00C3# else
		x"251A" when address_in = 16#00C4# else
		x"288D" when address_in = 16#00C5# else
		x"2B64" when address_in = 16#00C6# else
		x"2D93" when address_in = 16#00C7# else
		x"2F13" when address_in = 16#00C8# else
		x"2FDE" when address_in = 16#00C9# else
		x"2FF1" when address_in = 16#00CA# else
		x"2F4B" when address_in = 16#00CB# else
		x"2DEE" when address_in = 16#00CC# else
		x"2BE1" when address_in = 16#00CD# else
		x"292B" when address_in = 16#00CE# else
		x"25D7" when address_in = 16#00CF# else
		x"21F0" when address_in = 16#00D0# else
		x"1D87" when address_in = 16#00D1# else
		x"18AD" when address_in = 16#00D2# else
		x"1373" when address_in = 16#00D3# else
		x"0DEF" when address_in = 16#00D4# else
		x"0834" when address_in = 16#00D5# else
		x"025A" when address_in = 16#00D6# else
		x"FC79" when address_in = 16#00D7# else
		x"F6A3" when address_in = 16#00D8# else
		x"F0F2" when address_in = 16#00D9# else
		x"EB7B" when address_in = 16#00DA# else
		x"E652" when address_in = 16#00DB# else
		x"E18D" when address_in = 16#00DC# else
		x"DD3D" when address_in = 16#00DD# else
		x"D973" when address_in = 16#00DE# else
		x"D63D" when address_in = 16#00DF# else
		x"D3A8" when address_in = 16#00E0# else
		x"D1BE" when address_in = 16#00E1# else
		x"D085" when address_in = 16#00E2# else
		x"D004" when address_in = 16#00E3# else
		x"D03C" when address_in = 16#00E4# else
		x"D12B" when address_in = 16#00E5# else
		x"D2CF" when address_in = 16#00E6# else
		x"D521" when address_in = 16#00E7# else
		x"D817" when address_in = 16#00E8# else
		x"DBA8" when address_in = 16#00E9# else
		x"DFC4" when address_in = 16#00EA# else
		x"E45D" when address_in = 16#00EB# else
		x"E960" when address_in = 16#00EC# else
		x"EEBA" when address_in = 16#00ED# else
		x"F457" when address_in = 16#00EE# else
		x"FA20" when address_in = 16#00EF# else
		x"0000" when address_in = 16#00F0# else
		x"05E0" when address_in = 16#00F1# else
		x"0BA9" when address_in = 16#00F2# else
		x"1146" when address_in = 16#00F3# else
		x"16A0" when address_in = 16#00F4# else
		x"1BA3" when address_in = 16#00F5# else
		x"203C" when address_in = 16#00F6# else
		x"2458" when address_in = 16#00F7# else
		x"27E9" when address_in = 16#00F8# else
		x"2ADF" when address_in = 16#00F9# else
		x"2D31" when address_in = 16#00FA# else
		x"2ED5" when address_in = 16#00FB# else
		x"2FC4" when address_in = 16#00FC# else
		x"2FFC" when address_in = 16#00FD# else
		x"2F7B" when address_in = 16#00FE# else
		x"2E42" when address_in = 16#00FF# else
		x"2C58" when address_in = 16#0100# else
		x"29C3" when address_in = 16#0101# else
		x"268D" when address_in = 16#0102# else
		x"22C3" when address_in = 16#0103# else
		x"1E73" when address_in = 16#0104# else
		x"19AE" when address_in = 16#0105# else
		x"1485" when address_in = 16#0106# else
		x"0F0E" when address_in = 16#0107# else
		x"095D" when address_in = 16#0108# else
		x"0387" when address_in = 16#0109# else
		x"FDA6" when address_in = 16#010A# else
		x"F7CC" when address_in = 16#010B# else
		x"F211" when address_in = 16#010C# else
		x"EC8D" when address_in = 16#010D# else
		x"E753" when address_in = 16#010E# else
		x"E279" when address_in = 16#010F# else
		x"DE10" when address_in = 16#0110# else
		x"DA29" when address_in = 16#0111# else
		x"D6D5" when address_in = 16#0112# else
		x"D41F" when address_in = 16#0113# else
		x"D212" when address_in = 16#0114# else
		x"D0B5" when address_in = 16#0115# else
		x"D00F" when address_in = 16#0116# else
		x"D022" when address_in = 16#0117# else
		x"D0ED" when address_in = 16#0118# else
		x"D26D" when address_in = 16#0119# else
		x"D49C" when address_in = 16#011A# else
		x"D773" when address_in = 16#011B# else
		x"DAE6" when address_in = 16#011C# else
		x"DEE7" when address_in = 16#011D# else
		x"E369" when address_in = 16#011E# else
		x"E858" when address_in = 16#011F# else
		x"EDA2" when address_in = 16#0120# else
		x"F333" when address_in = 16#0121# else
		x"F8F5" when address_in = 16#0122# else
		x"FED3" when address_in = 16#0123# else
		x"04B4" when address_in = 16#0124# else
		x"0A84" when address_in = 16#0125# else
		x"102B" when address_in = 16#0126# else
		x"1594" when address_in = 16#0127# else
		x"1AAA" when address_in = 16#0128# else
		x"1F5A" when address_in = 16#0129# else
		x"2390" when address_in = 16#012A# else
		x"273E" when address_in = 16#012B# else
		x"2A55" when address_in = 16#012C# else
		x"2CC8" when address_in = 16#012D# else
		x"2E8F" when address_in = 16#012E# else
		x"2FA3" when address_in = 16#012F# else
		x"0000" when address_in = 16#0130# else
		x"00C9" when address_in = 16#0131# else
		x"0192" when address_in = 16#0132# else
		x"025B" when address_in = 16#0133# else
		x"0324" when address_in = 16#0134# else
		x"03ED" when address_in = 16#0135# else
		x"04B6" when address_in = 16#0136# else
		x"057E" when address_in = 16#0137# else
		x"0647" when address_in = 16#0138# else
		x"0710" when address_in = 16#0139# else
		x"07D9" when address_in = 16#013A# else
		x"08A1" when address_in = 16#013B# else
		x"096A" when address_in = 16#013C# else
		x"0A32" when address_in = 16#013D# else
		x"0AFB" when address_in = 16#013E# else
		x"0BC3" when address_in = 16#013F# else
		x"0C8B" when address_in = 16#0140# else
		x"0D53" when address_in = 16#0141# else
		x"0E1B" when address_in = 16#0142# else
		x"0EE3" when address_in = 16#0143# else
		x"0FAB" when address_in = 16#0144# else
		x"1072" when address_in = 16#0145# else
		x"1139" when address_in = 16#0146# else
		x"1200" when address_in = 16#0147# else
		x"12C7" when address_in = 16#0148# else
		x"138E" when address_in = 16#0149# else
		x"1455" when address_in = 16#014A# else
		x"151B" when address_in = 16#014B# else
		x"15E1" when address_in = 16#014C# else
		x"16A7" when address_in = 16#014D# else
		x"176D" when address_in = 16#014E# else
		x"1833" when address_in = 16#014F# else
		x"18F8" when address_in = 16#0150# else
		x"19BD" when address_in = 16#0151# else
		x"1A82" when address_in = 16#0152# else
		x"1B46" when address_in = 16#0153# else
		x"1C0B" when address_in = 16#0154# else
		x"1CCF" when address_in = 16#0155# else
		x"1D93" when address_in = 16#0156# else
		x"1E56" when address_in = 16#0157# else
		x"1F19" when address_in = 16#0158# else
		x"1FDC" when address_in = 16#0159# else
		x"209F" when address_in = 16#015A# else
		x"2161" when address_in = 16#015B# else
		x"2223" when address_in = 16#015C# else
		x"22E4" when address_in = 16#015D# else
		x"23A6" when address_in = 16#015E# else
		x"2467" when address_in = 16#015F# else
		x"2527" when address_in = 16#0160# else
		x"25E7" when address_in = 16#0161# else
		x"26A7" when address_in = 16#0162# else
		x"2767" when address_in = 16#0163# else
		x"2826" when address_in = 16#0164# else
		x"28E5" when address_in = 16#0165# else
		x"29A3" when address_in = 16#0166# else
		x"2A61" when address_in = 16#0167# else
		x"2B1E" when address_in = 16#0168# else
		x"2BDB" when address_in = 16#0169# else
		x"2C98" when address_in = 16#016A# else
		x"2D54" when address_in = 16#016B# else
		x"2E10" when address_in = 16#016C# else
		x"2ECC" when address_in = 16#016D# else
		x"2F86" when address_in = 16#016E# else
		x"3041" when address_in = 16#016F# else
		x"30FB" when address_in = 16#0170# else
		x"31B4" when address_in = 16#0171# else
		x"326D" when address_in = 16#0172# else
		x"3326" when address_in = 16#0173# else
		x"33DE" when address_in = 16#0174# else
		x"3496" when address_in = 16#0175# else
		x"354D" when address_in = 16#0176# else
		x"3603" when address_in = 16#0177# else
		x"36B9" when address_in = 16#0178# else
		x"376F" when address_in = 16#0179# else
		x"3824" when address_in = 16#017A# else
		x"38D8" when address_in = 16#017B# else
		x"398C" when address_in = 16#017C# else
		x"3A3F" when address_in = 16#017D# else
		x"3AF2" when address_in = 16#017E# else
		x"3BA4" when address_in = 16#017F# else
		x"3C56" when address_in = 16#0180# else
		x"3D07" when address_in = 16#0181# else
		x"3DB7" when address_in = 16#0182# else
		x"3E67" when address_in = 16#0183# else
		x"3F16" when address_in = 16#0184# else
		x"3FC5" when address_in = 16#0185# else
		x"4073" when address_in = 16#0186# else
		x"4120" when address_in = 16#0187# else
		x"41CD" when address_in = 16#0188# else
		x"4279" when address_in = 16#0189# else
		x"4325" when address_in = 16#018A# else
		x"43D0" when address_in = 16#018B# else
		x"447A" when address_in = 16#018C# else
		x"4523" when address_in = 16#018D# else
		x"45CC" when address_in = 16#018E# else
		x"4674" when address_in = 16#018F# else
		x"471C" when address_in = 16#0190# else
		x"47C3" when address_in = 16#0191# else
		x"4869" when address_in = 16#0192# else
		x"490E" when address_in = 16#0193# else
		x"49B3" when address_in = 16#0194# else
		x"4A57" when address_in = 16#0195# else
		x"4AFA" when address_in = 16#0196# else
		x"4B9D" when address_in = 16#0197# else
		x"4C3F" when address_in = 16#0198# else
		x"4CE0" when address_in = 16#0199# else
		x"4D80" when address_in = 16#019A# else
		x"4E20" when address_in = 16#019B# else
		x"4EBF" when address_in = 16#019C# else
		x"4F5D" when address_in = 16#019D# else
		x"4FFA" when address_in = 16#019E# else
		x"5097" when address_in = 16#019F# else
		x"5133" when address_in = 16#01A0# else
		x"51CE" when address_in = 16#01A1# else
		x"5268" when address_in = 16#01A2# else
		x"5301" when address_in = 16#01A3# else
		x"539A" when address_in = 16#01A4# else
		x"5432" when address_in = 16#01A5# else
		x"54C9" when address_in = 16#01A6# else
		x"555F" when address_in = 16#01A7# else
		x"55F4" when address_in = 16#01A8# else
		x"5689" when address_in = 16#01A9# else
		x"571D" when address_in = 16#01AA# else
		x"57B0" when address_in = 16#01AB# else
		x"5842" when address_in = 16#01AC# else
		x"58D3" when address_in = 16#01AD# else
		x"5963" when address_in = 16#01AE# else
		x"59F3" when address_in = 16#01AF# else
		x"5A81" when address_in = 16#01B0# else
		x"5B0F" when address_in = 16#01B1# else
		x"5B9C" when address_in = 16#01B2# else
		x"5C28" when address_in = 16#01B3# else
		x"5CB3" when address_in = 16#01B4# else
		x"5D3D" when address_in = 16#01B5# else
		x"5DC6" when address_in = 16#01B6# else
		x"5E4F" when address_in = 16#01B7# else
		x"5ED6" when address_in = 16#01B8# else
		x"5F5D" when address_in = 16#01B9# else
		x"5FE2" when address_in = 16#01BA# else
		x"6067" when address_in = 16#01BB# else
		x"60EB" when address_in = 16#01BC# else
		x"616E" when address_in = 16#01BD# else
		x"61F0" when address_in = 16#01BE# else
		x"6271" when address_in = 16#01BF# else
		x"62F1" when address_in = 16#01C0# else
		x"6370" when address_in = 16#01C1# else
		x"63EE" when address_in = 16#01C2# else
		x"646B" when address_in = 16#01C3# else
		x"64E7" when address_in = 16#01C4# else
		x"6562" when address_in = 16#01C5# else
		x"65DD" when address_in = 16#01C6# else
		x"6656" when address_in = 16#01C7# else
		x"66CE" when address_in = 16#01C8# else
		x"6745" when address_in = 16#01C9# else
		x"67BC" when address_in = 16#01CA# else
		x"6831" when address_in = 16#01CB# else
		x"68A5" when address_in = 16#01CC# else
		x"6919" when address_in = 16#01CD# else
		x"698B" when address_in = 16#01CE# else
		x"69FC" when address_in = 16#01CF# else
		x"6A6C" when address_in = 16#01D0# else
		x"6ADB" when address_in = 16#01D1# else
		x"6B4A" when address_in = 16#01D2# else
		x"6BB7" when address_in = 16#01D3# else
		x"6C23" when address_in = 16#01D4# else
		x"6C8E" when address_in = 16#01D5# else
		x"6CF8" when address_in = 16#01D6# else
		x"6D61" when address_in = 16#01D7# else
		x"6DC9" when address_in = 16#01D8# else
		x"6E30" when address_in = 16#01D9# else
		x"6E95" when address_in = 16#01DA# else
		x"6EFA" when address_in = 16#01DB# else
		x"6F5E" when address_in = 16#01DC# else
		x"6FC0" when address_in = 16#01DD# else
		x"7022" when address_in = 16#01DE# else
		x"7082" when address_in = 16#01DF# else
		x"70E1" when address_in = 16#01E0# else
		x"7140" when address_in = 16#01E1# else
		x"719D" when address_in = 16#01E2# else
		x"71F9" when address_in = 16#01E3# else
		x"7254" when address_in = 16#01E4# else
		x"72AE" when address_in = 16#01E5# else
		x"7306" when address_in = 16#01E6# else
		x"735E" when address_in = 16#01E7# else
		x"73B5" when address_in = 16#01E8# else
		x"740A" when address_in = 16#01E9# else
		x"745E" when address_in = 16#01EA# else
		x"74B1" when address_in = 16#01EB# else
		x"7503" when address_in = 16#01EC# else
		x"7554" when address_in = 16#01ED# else
		x"75A4" when address_in = 16#01EE# else
		x"75F3" when address_in = 16#01EF# else
		x"7640" when address_in = 16#01F0# else
		x"768D" when address_in = 16#01F1# else
		x"76D8" when address_in = 16#01F2# else
		x"7722" when address_in = 16#01F3# else
		x"776B" when address_in = 16#01F4# else
		x"77B3" when address_in = 16#01F5# else
		x"77F9" when address_in = 16#01F6# else
		x"783F" when address_in = 16#01F7# else
		x"7883" when address_in = 16#01F8# else
		x"78C6" when address_in = 16#01F9# else
		x"7908" when address_in = 16#01FA# else
		x"7949" when address_in = 16#01FB# else
		x"7989" when address_in = 16#01FC# else
		x"79C7" when address_in = 16#01FD# else
		x"7A04" when address_in = 16#01FE# else
		x"7A41" when address_in = 16#01FF# else
		x"7A7C" when address_in = 16#0200# else
		x"7AB5" when address_in = 16#0201# else
		x"7AEE" when address_in = 16#0202# else
		x"7B25" when address_in = 16#0203# else
		x"7B5C" when address_in = 16#0204# else
		x"7B91" when address_in = 16#0205# else
		x"7BC4" when address_in = 16#0206# else
		x"7BF7" when address_in = 16#0207# else
		x"7C29" when address_in = 16#0208# else
		x"7C59" when address_in = 16#0209# else
		x"7C88" when address_in = 16#020A# else
		x"7CB6" when address_in = 16#020B# else
		x"7CE2" when address_in = 16#020C# else
		x"7D0E" when address_in = 16#020D# else
		x"7D38" when address_in = 16#020E# else
		x"7D61" when address_in = 16#020F# else
		x"7D89" when address_in = 16#0210# else
		x"7DB0" when address_in = 16#0211# else
		x"7DD5" when address_in = 16#0212# else
		x"7DF9" when address_in = 16#0213# else
		x"7E1C" when address_in = 16#0214# else
		x"7E3E" when address_in = 16#0215# else
		x"7E5E" when address_in = 16#0216# else
		x"7E7E" when address_in = 16#0217# else
		x"7E9C" when address_in = 16#0218# else
		x"7EB9" when address_in = 16#0219# else
		x"7ED4" when address_in = 16#021A# else
		x"7EEF" when address_in = 16#021B# else
		x"7F08" when address_in = 16#021C# else
		x"7F20" when address_in = 16#021D# else
		x"7F37" when address_in = 16#021E# else
		x"7F4C" when address_in = 16#021F# else
		x"7F61" when address_in = 16#0220# else
		x"7F74" when address_in = 16#0221# else
		x"7F86" when address_in = 16#0222# else
		x"7F96" when address_in = 16#0223# else
		x"7FA6" when address_in = 16#0224# else
		x"7FB4" when address_in = 16#0225# else
		x"7FC1" when address_in = 16#0226# else
		x"7FCD" when address_in = 16#0227# else
		x"7FD7" when address_in = 16#0228# else
		x"7FE0" when address_in = 16#0229# else
		x"7FE8" when address_in = 16#022A# else
		x"7FEF" when address_in = 16#022B# else
		x"7FF5" when address_in = 16#022C# else
		x"7FF9" when address_in = 16#022D# else
		x"7FFC" when address_in = 16#022E# else
		x"7FFE" when address_in = 16#022F# else
		x"7FFF" when address_in = 16#0230# else
		x"7FFE" when address_in = 16#0231# else
		x"7FFC" when address_in = 16#0232# else
		x"7FF9" when address_in = 16#0233# else
		x"7FF5" when address_in = 16#0234# else
		x"7FEF" when address_in = 16#0235# else
		x"7FE8" when address_in = 16#0236# else
		x"7FE0" when address_in = 16#0237# else
		x"7FD7" when address_in = 16#0238# else
		x"7FCD" when address_in = 16#0239# else
		x"7FC1" when address_in = 16#023A# else
		x"7FB4" when address_in = 16#023B# else
		x"7FA6" when address_in = 16#023C# else
		x"7F96" when address_in = 16#023D# else
		x"7F86" when address_in = 16#023E# else
		x"7F74" when address_in = 16#023F# else
		x"7F61" when address_in = 16#0240# else
		x"7F4C" when address_in = 16#0241# else
		x"7F37" when address_in = 16#0242# else
		x"7F20" when address_in = 16#0243# else
		x"7F08" when address_in = 16#0244# else
		x"7EEF" when address_in = 16#0245# else
		x"7ED4" when address_in = 16#0246# else
		x"7EB9" when address_in = 16#0247# else
		x"7E9C" when address_in = 16#0248# else
		x"7E7E" when address_in = 16#0249# else
		x"7E5E" when address_in = 16#024A# else
		x"7E3E" when address_in = 16#024B# else
		x"7E1C" when address_in = 16#024C# else
		x"7DF9" when address_in = 16#024D# else
		x"7DD5" when address_in = 16#024E# else
		x"7DB0" when address_in = 16#024F# else
		x"7D89" when address_in = 16#0250# else
		x"7D61" when address_in = 16#0251# else
		x"7D38" when address_in = 16#0252# else
		x"7D0E" when address_in = 16#0253# else
		x"7CE2" when address_in = 16#0254# else
		x"7CB6" when address_in = 16#0255# else
		x"7C88" when address_in = 16#0256# else
		x"7C59" when address_in = 16#0257# else
		x"7C29" when address_in = 16#0258# else
		x"7BF7" when address_in = 16#0259# else
		x"7BC4" when address_in = 16#025A# else
		x"7B91" when address_in = 16#025B# else
		x"7B5C" when address_in = 16#025C# else
		x"7B25" when address_in = 16#025D# else
		x"7AEE" when address_in = 16#025E# else
		x"7AB5" when address_in = 16#025F# else
		x"7A7C" when address_in = 16#0260# else
		x"7A41" when address_in = 16#0261# else
		x"7A04" when address_in = 16#0262# else
		x"79C7" when address_in = 16#0263# else
		x"7989" when address_in = 16#0264# else
		x"7949" when address_in = 16#0265# else
		x"7908" when address_in = 16#0266# else
		x"78C6" when address_in = 16#0267# else
		x"7883" when address_in = 16#0268# else
		x"783F" when address_in = 16#0269# else
		x"77F9" when address_in = 16#026A# else
		x"77B3" when address_in = 16#026B# else
		x"776B" when address_in = 16#026C# else
		x"7722" when address_in = 16#026D# else
		x"76D8" when address_in = 16#026E# else
		x"768D" when address_in = 16#026F# else
		x"7640" when address_in = 16#0270# else
		x"75F3" when address_in = 16#0271# else
		x"75A4" when address_in = 16#0272# else
		x"7554" when address_in = 16#0273# else
		x"7503" when address_in = 16#0274# else
		x"74B1" when address_in = 16#0275# else
		x"745E" when address_in = 16#0276# else
		x"740A" when address_in = 16#0277# else
		x"73B5" when address_in = 16#0278# else
		x"735E" when address_in = 16#0279# else
		x"7306" when address_in = 16#027A# else
		x"72AE" when address_in = 16#027B# else
		x"7254" when address_in = 16#027C# else
		x"71F9" when address_in = 16#027D# else
		x"719D" when address_in = 16#027E# else
		x"7140" when address_in = 16#027F# else
		x"70E1" when address_in = 16#0280# else
		x"7082" when address_in = 16#0281# else
		x"7022" when address_in = 16#0282# else
		x"6FC0" when address_in = 16#0283# else
		x"6F5E" when address_in = 16#0284# else
		x"6EFA" when address_in = 16#0285# else
		x"6E95" when address_in = 16#0286# else
		x"6E30" when address_in = 16#0287# else
		x"6DC9" when address_in = 16#0288# else
		x"6D61" when address_in = 16#0289# else
		x"6CF8" when address_in = 16#028A# else
		x"6C8E" when address_in = 16#028B# else
		x"6C23" when address_in = 16#028C# else
		x"6BB7" when address_in = 16#028D# else
		x"6B4A" when address_in = 16#028E# else
		x"6ADB" when address_in = 16#028F# else
		x"6A6C" when address_in = 16#0290# else
		x"69FC" when address_in = 16#0291# else
		x"698B" when address_in = 16#0292# else
		x"6919" when address_in = 16#0293# else
		x"68A5" when address_in = 16#0294# else
		x"6831" when address_in = 16#0295# else
		x"67BC" when address_in = 16#0296# else
		x"6745" when address_in = 16#0297# else
		x"66CE" when address_in = 16#0298# else
		x"6656" when address_in = 16#0299# else
		x"65DD" when address_in = 16#029A# else
		x"6562" when address_in = 16#029B# else
		x"64E7" when address_in = 16#029C# else
		x"646B" when address_in = 16#029D# else
		x"63EE" when address_in = 16#029E# else
		x"6370" when address_in = 16#029F# else
		x"62F1" when address_in = 16#02A0# else
		x"6271" when address_in = 16#02A1# else
		x"61F0" when address_in = 16#02A2# else
		x"616E" when address_in = 16#02A3# else
		x"60EB" when address_in = 16#02A4# else
		x"6067" when address_in = 16#02A5# else
		x"5FE2" when address_in = 16#02A6# else
		x"5F5D" when address_in = 16#02A7# else
		x"5ED6" when address_in = 16#02A8# else
		x"5E4F" when address_in = 16#02A9# else
		x"5DC6" when address_in = 16#02AA# else
		x"5D3D" when address_in = 16#02AB# else
		x"5CB3" when address_in = 16#02AC# else
		x"5C28" when address_in = 16#02AD# else
		x"5B9C" when address_in = 16#02AE# else
		x"5B0F" when address_in = 16#02AF# else
		x"5A81" when address_in = 16#02B0# else
		x"59F3" when address_in = 16#02B1# else
		x"5963" when address_in = 16#02B2# else
		x"58D3" when address_in = 16#02B3# else
		x"5842" when address_in = 16#02B4# else
		x"57B0" when address_in = 16#02B5# else
		x"571D" when address_in = 16#02B6# else
		x"5689" when address_in = 16#02B7# else
		x"55F4" when address_in = 16#02B8# else
		x"555F" when address_in = 16#02B9# else
		x"54C9" when address_in = 16#02BA# else
		x"5432" when address_in = 16#02BB# else
		x"539A" when address_in = 16#02BC# else
		x"5301" when address_in = 16#02BD# else
		x"5268" when address_in = 16#02BE# else
		x"51CE" when address_in = 16#02BF# else
		x"5133" when address_in = 16#02C0# else
		x"5097" when address_in = 16#02C1# else
		x"4FFA" when address_in = 16#02C2# else
		x"4F5D" when address_in = 16#02C3# else
		x"4EBF" when address_in = 16#02C4# else
		x"4E20" when address_in = 16#02C5# else
		x"4D80" when address_in = 16#02C6# else
		x"4CE0" when address_in = 16#02C7# else
		x"4C3F" when address_in = 16#02C8# else
		x"4B9D" when address_in = 16#02C9# else
		x"4AFA" when address_in = 16#02CA# else
		x"4A57" when address_in = 16#02CB# else
		x"49B3" when address_in = 16#02CC# else
		x"490E" when address_in = 16#02CD# else
		x"4869" when address_in = 16#02CE# else
		x"47C3" when address_in = 16#02CF# else
		x"471C" when address_in = 16#02D0# else
		x"4674" when address_in = 16#02D1# else
		x"45CC" when address_in = 16#02D2# else
		x"4523" when address_in = 16#02D3# else
		x"447A" when address_in = 16#02D4# else
		x"43D0" when address_in = 16#02D5# else
		x"4325" when address_in = 16#02D6# else
		x"4279" when address_in = 16#02D7# else
		x"41CD" when address_in = 16#02D8# else
		x"4120" when address_in = 16#02D9# else
		x"4073" when address_in = 16#02DA# else
		x"3FC5" when address_in = 16#02DB# else
		x"3F16" when address_in = 16#02DC# else
		x"3E67" when address_in = 16#02DD# else
		x"3DB7" when address_in = 16#02DE# else
		x"3D07" when address_in = 16#02DF# else
		x"3C56" when address_in = 16#02E0# else
		x"3BA4" when address_in = 16#02E1# else
		x"3AF2" when address_in = 16#02E2# else
		x"3A3F" when address_in = 16#02E3# else
		x"398C" when address_in = 16#02E4# else
		x"38D8" when address_in = 16#02E5# else
		x"3824" when address_in = 16#02E6# else
		x"376F" when address_in = 16#02E7# else
		x"36B9" when address_in = 16#02E8# else
		x"3603" when address_in = 16#02E9# else
		x"354D" when address_in = 16#02EA# else
		x"3496" when address_in = 16#02EB# else
		x"33DE" when address_in = 16#02EC# else
		x"3326" when address_in = 16#02ED# else
		x"326D" when address_in = 16#02EE# else
		x"31B4" when address_in = 16#02EF# else
		x"30FB" when address_in = 16#02F0# else
		x"3041" when address_in = 16#02F1# else
		x"2F86" when address_in = 16#02F2# else
		x"2ECC" when address_in = 16#02F3# else
		x"2E10" when address_in = 16#02F4# else
		x"2D54" when address_in = 16#02F5# else
		x"2C98" when address_in = 16#02F6# else
		x"2BDB" when address_in = 16#02F7# else
		x"2B1E" when address_in = 16#02F8# else
		x"2A61" when address_in = 16#02F9# else
		x"29A3" when address_in = 16#02FA# else
		x"28E5" when address_in = 16#02FB# else
		x"2826" when address_in = 16#02FC# else
		x"2767" when address_in = 16#02FD# else
		x"26A7" when address_in = 16#02FE# else
		x"25E7" when address_in = 16#02FF# else
		x"2527" when address_in = 16#0300# else
		x"2467" when address_in = 16#0301# else
		x"23A6" when address_in = 16#0302# else
		x"22E4" when address_in = 16#0303# else
		x"2223" when address_in = 16#0304# else
		x"2161" when address_in = 16#0305# else
		x"209F" when address_in = 16#0306# else
		x"1FDC" when address_in = 16#0307# else
		x"1F19" when address_in = 16#0308# else
		x"1E56" when address_in = 16#0309# else
		x"1D93" when address_in = 16#030A# else
		x"1CCF" when address_in = 16#030B# else
		x"1C0B" when address_in = 16#030C# else
		x"1B46" when address_in = 16#030D# else
		x"1A82" when address_in = 16#030E# else
		x"19BD" when address_in = 16#030F# else
		x"18F8" when address_in = 16#0310# else
		x"1833" when address_in = 16#0311# else
		x"176D" when address_in = 16#0312# else
		x"16A7" when address_in = 16#0313# else
		x"15E1" when address_in = 16#0314# else
		x"151B" when address_in = 16#0315# else
		x"1455" when address_in = 16#0316# else
		x"138E" when address_in = 16#0317# else
		x"12C7" when address_in = 16#0318# else
		x"1200" when address_in = 16#0319# else
		x"1139" when address_in = 16#031A# else
		x"1072" when address_in = 16#031B# else
		x"0FAB" when address_in = 16#031C# else
		x"0EE3" when address_in = 16#031D# else
		x"0E1B" when address_in = 16#031E# else
		x"0D53" when address_in = 16#031F# else
		x"0C8B" when address_in = 16#0320# else
		x"0BC3" when address_in = 16#0321# else
		x"0AFB" when address_in = 16#0322# else
		x"0A32" when address_in = 16#0323# else
		x"096A" when address_in = 16#0324# else
		x"08A1" when address_in = 16#0325# else
		x"07D9" when address_in = 16#0326# else
		x"0710" when address_in = 16#0327# else
		x"0647" when address_in = 16#0328# else
		x"057E" when address_in = 16#0329# else
		x"04B6" when address_in = 16#032A# else
		x"03ED" when address_in = 16#032B# else
		x"0324" when address_in = 16#032C# else
		x"025B" when address_in = 16#032D# else
		x"0192" when address_in = 16#032E# else
		x"00C9" when address_in = 16#032F# else
		x"0000" when address_in = 16#0330# else
		x"FF37" when address_in = 16#0331# else
		x"FE6E" when address_in = 16#0332# else
		x"FDA5" when address_in = 16#0333# else
		x"FCDC" when address_in = 16#0334# else
		x"FC13" when address_in = 16#0335# else
		x"FB4A" when address_in = 16#0336# else
		x"FA82" when address_in = 16#0337# else
		x"F9B9" when address_in = 16#0338# else
		x"F8F0" when address_in = 16#0339# else
		x"F827" when address_in = 16#033A# else
		x"F75F" when address_in = 16#033B# else
		x"F696" when address_in = 16#033C# else
		x"F5CE" when address_in = 16#033D# else
		x"F505" when address_in = 16#033E# else
		x"F43D" when address_in = 16#033F# else
		x"F375" when address_in = 16#0340# else
		x"F2AD" when address_in = 16#0341# else
		x"F1E5" when address_in = 16#0342# else
		x"F11D" when address_in = 16#0343# else
		x"F055" when address_in = 16#0344# else
		x"EF8E" when address_in = 16#0345# else
		x"EEC7" when address_in = 16#0346# else
		x"EE00" when address_in = 16#0347# else
		x"ED39" when address_in = 16#0348# else
		x"EC72" when address_in = 16#0349# else
		x"EBAB" when address_in = 16#034A# else
		x"EAE5" when address_in = 16#034B# else
		x"EA1F" when address_in = 16#034C# else
		x"E959" when address_in = 16#034D# else
		x"E893" when address_in = 16#034E# else
		x"E7CD" when address_in = 16#034F# else
		x"E708" when address_in = 16#0350# else
		x"E643" when address_in = 16#0351# else
		x"E57E" when address_in = 16#0352# else
		x"E4BA" when address_in = 16#0353# else
		x"E3F5" when address_in = 16#0354# else
		x"E331" when address_in = 16#0355# else
		x"E26D" when address_in = 16#0356# else
		x"E1AA" when address_in = 16#0357# else
		x"E0E7" when address_in = 16#0358# else
		x"E024" when address_in = 16#0359# else
		x"DF61" when address_in = 16#035A# else
		x"DE9F" when address_in = 16#035B# else
		x"DDDD" when address_in = 16#035C# else
		x"DD1C" when address_in = 16#035D# else
		x"DC5A" when address_in = 16#035E# else
		x"DB99" when address_in = 16#035F# else
		x"DAD9" when address_in = 16#0360# else
		x"DA19" when address_in = 16#0361# else
		x"D959" when address_in = 16#0362# else
		x"D899" when address_in = 16#0363# else
		x"D7DA" when address_in = 16#0364# else
		x"D71B" when address_in = 16#0365# else
		x"D65D" when address_in = 16#0366# else
		x"D59F" when address_in = 16#0367# else
		x"D4E2" when address_in = 16#0368# else
		x"D425" when address_in = 16#0369# else
		x"D368" when address_in = 16#036A# else
		x"D2AC" when address_in = 16#036B# else
		x"D1F0" when address_in = 16#036C# else
		x"D134" when address_in = 16#036D# else
		x"D07A" when address_in = 16#036E# else
		x"CFBF" when address_in = 16#036F# else
		x"CF05" when address_in = 16#0370# else
		x"CE4C" when address_in = 16#0371# else
		x"CD93" when address_in = 16#0372# else
		x"CCDA" when address_in = 16#0373# else
		x"CC22" when address_in = 16#0374# else
		x"CB6A" when address_in = 16#0375# else
		x"CAB3" when address_in = 16#0376# else
		x"C9FD" when address_in = 16#0377# else
		x"C947" when address_in = 16#0378# else
		x"C891" when address_in = 16#0379# else
		x"C7DC" when address_in = 16#037A# else
		x"C728" when address_in = 16#037B# else
		x"C674" when address_in = 16#037C# else
		x"C5C1" when address_in = 16#037D# else
		x"C50E" when address_in = 16#037E# else
		x"C45C" when address_in = 16#037F# else
		x"C3AA" when address_in = 16#0380# else
		x"C2F9" when address_in = 16#0381# else
		x"C249" when address_in = 16#0382# else
		x"C199" when address_in = 16#0383# else
		x"C0EA" when address_in = 16#0384# else
		x"C03B" when address_in = 16#0385# else
		x"BF8D" when address_in = 16#0386# else
		x"BEE0" when address_in = 16#0387# else
		x"BE33" when address_in = 16#0388# else
		x"BD87" when address_in = 16#0389# else
		x"BCDB" when address_in = 16#038A# else
		x"BC30" when address_in = 16#038B# else
		x"BB86" when address_in = 16#038C# else
		x"BADD" when address_in = 16#038D# else
		x"BA34" when address_in = 16#038E# else
		x"B98C" when address_in = 16#038F# else
		x"B8E4" when address_in = 16#0390# else
		x"B83D" when address_in = 16#0391# else
		x"B797" when address_in = 16#0392# else
		x"B6F2" when address_in = 16#0393# else
		x"B64D" when address_in = 16#0394# else
		x"B5A9" when address_in = 16#0395# else
		x"B506" when address_in = 16#0396# else
		x"B463" when address_in = 16#0397# else
		x"B3C1" when address_in = 16#0398# else
		x"B320" when address_in = 16#0399# else
		x"B280" when address_in = 16#039A# else
		x"B1E0" when address_in = 16#039B# else
		x"B141" when address_in = 16#039C# else
		x"B0A3" when address_in = 16#039D# else
		x"B006" when address_in = 16#039E# else
		x"AF69" when address_in = 16#039F# else
		x"AECD" when address_in = 16#03A0# else
		x"AE32" when address_in = 16#03A1# else
		x"AD98" when address_in = 16#03A2# else
		x"ACFF" when address_in = 16#03A3# else
		x"AC66" when address_in = 16#03A4# else
		x"ABCE" when address_in = 16#03A5# else
		x"AB37" when address_in = 16#03A6# else
		x"AAA1" when address_in = 16#03A7# else
		x"AA0C" when address_in = 16#03A8# else
		x"A977" when address_in = 16#03A9# else
		x"A8E3" when address_in = 16#03AA# else
		x"A850" when address_in = 16#03AB# else
		x"A7BE" when address_in = 16#03AC# else
		x"A72D" when address_in = 16#03AD# else
		x"A69D" when address_in = 16#03AE# else
		x"A60D" when address_in = 16#03AF# else
		x"A57F" when address_in = 16#03B0# else
		x"A4F1" when address_in = 16#03B1# else
		x"A464" when address_in = 16#03B2# else
		x"A3D8" when address_in = 16#03B3# else
		x"A34D" when address_in = 16#03B4# else
		x"A2C3" when address_in = 16#03B5# else
		x"A23A" when address_in = 16#03B6# else
		x"A1B1" when address_in = 16#03B7# else
		x"A12A" when address_in = 16#03B8# else
		x"A0A3" when address_in = 16#03B9# else
		x"A01E" when address_in = 16#03BA# else
		x"9F99" when address_in = 16#03BB# else
		x"9F15" when address_in = 16#03BC# else
		x"9E92" when address_in = 16#03BD# else
		x"9E10" when address_in = 16#03BE# else
		x"9D8F" when address_in = 16#03BF# else
		x"9D0F" when address_in = 16#03C0# else
		x"9C90" when address_in = 16#03C1# else
		x"9C12" when address_in = 16#03C2# else
		x"9B95" when address_in = 16#03C3# else
		x"9B19" when address_in = 16#03C4# else
		x"9A9E" when address_in = 16#03C5# else
		x"9A23" when address_in = 16#03C6# else
		x"99AA" when address_in = 16#03C7# else
		x"9932" when address_in = 16#03C8# else
		x"98BB" when address_in = 16#03C9# else
		x"9844" when address_in = 16#03CA# else
		x"97CF" when address_in = 16#03CB# else
		x"975B" when address_in = 16#03CC# else
		x"96E7" when address_in = 16#03CD# else
		x"9675" when address_in = 16#03CE# else
		x"9604" when address_in = 16#03CF# else
		x"9594" when address_in = 16#03D0# else
		x"9525" when address_in = 16#03D1# else
		x"94B6" when address_in = 16#03D2# else
		x"9449" when address_in = 16#03D3# else
		x"93DD" when address_in = 16#03D4# else
		x"9372" when address_in = 16#03D5# else
		x"9308" when address_in = 16#03D6# else
		x"929F" when address_in = 16#03D7# else
		x"9237" when address_in = 16#03D8# else
		x"91D0" when address_in = 16#03D9# else
		x"916B" when address_in = 16#03DA# else
		x"9106" when address_in = 16#03DB# else
		x"90A2" when address_in = 16#03DC# else
		x"9040" when address_in = 16#03DD# else
		x"8FDE" when address_in = 16#03DE# else
		x"8F7E" when address_in = 16#03DF# else
		x"8F1F" when address_in = 16#03E0# else
		x"8EC0" when address_in = 16#03E1# else
		x"8E63" when address_in = 16#03E2# else
		x"8E07" when address_in = 16#03E3# else
		x"8DAC" when address_in = 16#03E4# else
		x"8D52" when address_in = 16#03E5# else
		x"8CFA" when address_in = 16#03E6# else
		x"8CA2" when address_in = 16#03E7# else
		x"8C4B" when address_in = 16#03E8# else
		x"8BF6" when address_in = 16#03E9# else
		x"8BA2" when address_in = 16#03EA# else
		x"8B4F" when address_in = 16#03EB# else
		x"8AFD" when address_in = 16#03EC# else
		x"8AAC" when address_in = 16#03ED# else
		x"8A5C" when address_in = 16#03EE# else
		x"8A0D" when address_in = 16#03EF# else
		x"89C0" when address_in = 16#03F0# else
		x"8973" when address_in = 16#03F1# else
		x"8928" when address_in = 16#03F2# else
		x"88DE" when address_in = 16#03F3# else
		x"8895" when address_in = 16#03F4# else
		x"884D" when address_in = 16#03F5# else
		x"8807" when address_in = 16#03F6# else
		x"87C1" when address_in = 16#03F7# else
		x"877D" when address_in = 16#03F8# else
		x"873A" when address_in = 16#03F9# else
		x"86F8" when address_in = 16#03FA# else
		x"86B7" when address_in = 16#03FB# else
		x"8677" when address_in = 16#03FC# else
		x"8639" when address_in = 16#03FD# else
		x"85FC" when address_in = 16#03FE# else
		x"85BF" when address_in = 16#03FF# else
		x"8584" when address_in = 16#0400# else
		x"854B" when address_in = 16#0401# else
		x"8512" when address_in = 16#0402# else
		x"84DB" when address_in = 16#0403# else
		x"84A4" when address_in = 16#0404# else
		x"846F" when address_in = 16#0405# else
		x"843C" when address_in = 16#0406# else
		x"8409" when address_in = 16#0407# else
		x"83D7" when address_in = 16#0408# else
		x"83A7" when address_in = 16#0409# else
		x"8378" when address_in = 16#040A# else
		x"834A" when address_in = 16#040B# else
		x"831E" when address_in = 16#040C# else
		x"82F2" when address_in = 16#040D# else
		x"82C8" when address_in = 16#040E# else
		x"829F" when address_in = 16#040F# else
		x"8277" when address_in = 16#0410# else
		x"8250" when address_in = 16#0411# else
		x"822B" when address_in = 16#0412# else
		x"8207" when address_in = 16#0413# else
		x"81E4" when address_in = 16#0414# else
		x"81C2" when address_in = 16#0415# else
		x"81A2" when address_in = 16#0416# else
		x"8182" when address_in = 16#0417# else
		x"8164" when address_in = 16#0418# else
		x"8147" when address_in = 16#0419# else
		x"812C" when address_in = 16#041A# else
		x"8111" when address_in = 16#041B# else
		x"80F8" when address_in = 16#041C# else
		x"80E0" when address_in = 16#041D# else
		x"80C9" when address_in = 16#041E# else
		x"80B4" when address_in = 16#041F# else
		x"809F" when address_in = 16#0420# else
		x"808C" when address_in = 16#0421# else
		x"807A" when address_in = 16#0422# else
		x"806A" when address_in = 16#0423# else
		x"805A" when address_in = 16#0424# else
		x"804C" when address_in = 16#0425# else
		x"803F" when address_in = 16#0426# else
		x"8033" when address_in = 16#0427# else
		x"8029" when address_in = 16#0428# else
		x"8020" when address_in = 16#0429# else
		x"8018" when address_in = 16#042A# else
		x"8011" when address_in = 16#042B# else
		x"800B" when address_in = 16#042C# else
		x"8007" when address_in = 16#042D# else
		x"8004" when address_in = 16#042E# else
		x"8002" when address_in = 16#042F# else
		x"2411" when address_in = 16#0430# else
		x"BE1F" when address_in = 16#0431# else
		x"EFCF" when address_in = 16#0432# else
		x"E0DF" when address_in = 16#0433# else
		x"BFDE" when address_in = 16#0434# else
		x"BFCD" when address_in = 16#0435# else
		x"E011" when address_in = 16#0436# else
		x"E6A0" when address_in = 16#0437# else
		x"E0B0" when address_in = 16#0438# else
		x"E2E8" when address_in = 16#0439# else
		x"E1F6" when address_in = 16#043A# else
		x"EF0F" when address_in = 16#043B# else
		x"9503" when address_in = 16#043C# else
		x"BF0B" when address_in = 16#043D# else
		x"C004" when address_in = 16#043E# else
		x"95D8" when address_in = 16#043F# else
		x"920D" when address_in = 16#0440# else
		x"9631" when address_in = 16#0441# else
		x"F3C8" when address_in = 16#0442# else
		x"36A0" when address_in = 16#0443# else
		x"07B1" when address_in = 16#0444# else
		x"F7C9" when address_in = 16#0445# else
		x"E011" when address_in = 16#0446# else
		x"E6A0" when address_in = 16#0447# else
		x"E0B1" when address_in = 16#0448# else
		x"C001" when address_in = 16#0449# else
		x"921D" when address_in = 16#044A# else
		x"36A6" when address_in = 16#044B# else
		x"07B1" when address_in = 16#044C# else
		x"F7E1" when address_in = 16#044D# else
		x"940C" when address_in = 16#044E# else
		x"0458" when address_in = 16#044F# else
		x"940C" when address_in = 16#0450# else
		x"0000" when address_in = 16#0451# else
		x"FF97" when address_in = 16#0452# else
		x"C003" when address_in = 16#0453# else
		x"9590" when address_in = 16#0454# else
		x"9581" when address_in = 16#0455# else
		x"4F9F" when address_in = 16#0456# else
		x"9508" when address_in = 16#0457# else
		x"EFCF" when address_in = 16#0458# else
		x"E0DF" when address_in = 16#0459# else
		x"BFDE" when address_in = 16#045A# else
		x"BFCD" when address_in = 16#045B# else
		x"E688" when address_in = 16#045C# else
		x"B983" when address_in = 16#045D# else
		x"E089" when address_in = 16#045E# else
		x"B982" when address_in = 16#045F# else
		x"940E" when address_in = 16#0460# else
		x"0728" when address_in = 16#0461# else
		x"940E" when address_in = 16#0462# else
		x"1000" when address_in = 16#0463# else
		x"CFFF" when address_in = 16#0464# else
		x"928F" when address_in = 16#0465# else
		x"929F" when address_in = 16#0466# else
		x"92AF" when address_in = 16#0467# else
		x"92BF" when address_in = 16#0468# else
		x"92CF" when address_in = 16#0469# else
		x"92DF" when address_in = 16#046A# else
		x"92EF" when address_in = 16#046B# else
		x"92FF" when address_in = 16#046C# else
		x"930F" when address_in = 16#046D# else
		x"931F" when address_in = 16#046E# else
		x"93CF" when address_in = 16#046F# else
		x"93DF" when address_in = 16#0470# else
		x"B184" when address_in = 16#0471# else
		x"2799" when address_in = 16#0472# else
		x"718E" when address_in = 16#0473# else
		x"7090" when address_in = 16#0474# else
		x"9595" when address_in = 16#0475# else
		x"9587" when address_in = 16#0476# else
		x"9595" when address_in = 16#0477# else
		x"9587" when address_in = 16#0478# else
		x"2F68" when address_in = 16#0479# else
		x"E080" when address_in = 16#047A# else
		x"E092" when address_in = 16#047B# else
		x"940E" when address_in = 16#047C# else
		x"1380" when address_in = 16#047D# else
		x"2EE8" when address_in = 16#047E# else
		x"2EF9" when address_in = 16#047F# else
		x"B184" when address_in = 16#0480# else
		x"2799" when address_in = 16#0481# else
		x"718E" when address_in = 16#0482# else
		x"7090" when address_in = 16#0483# else
		x"9595" when address_in = 16#0484# else
		x"9587" when address_in = 16#0485# else
		x"9595" when address_in = 16#0486# else
		x"9587" when address_in = 16#0487# else
		x"2F68" when address_in = 16#0488# else
		x"E080" when address_in = 16#0489# else
		x"E092" when address_in = 16#048A# else
		x"940E" when address_in = 16#048B# else
		x"1380" when address_in = 16#048C# else
		x"2F08" when address_in = 16#048D# else
		x"2F19" when address_in = 16#048E# else
		x"B184" when address_in = 16#048F# else
		x"2799" when address_in = 16#0490# else
		x"718E" when address_in = 16#0491# else
		x"7090" when address_in = 16#0492# else
		x"9595" when address_in = 16#0493# else
		x"9587" when address_in = 16#0494# else
		x"9595" when address_in = 16#0495# else
		x"9587" when address_in = 16#0496# else
		x"2F68" when address_in = 16#0497# else
		x"E082" when address_in = 16#0498# else
		x"E090" when address_in = 16#0499# else
		x"940E" when address_in = 16#049A# else
		x"1380" when address_in = 16#049B# else
		x"2EC8" when address_in = 16#049C# else
		x"2ED9" when address_in = 16#049D# else
		x"EF8F" when address_in = 16#049E# else
		x"BB8A" when address_in = 16#049F# else
		x"BA1B" when address_in = 16#04A0# else
		x"E0C0" when address_in = 16#04A1# else
		x"E0D0" when address_in = 16#04A2# else
		x"E040" when address_in = 16#04A3# else
		x"E051" when address_in = 16#04A4# else
		x"2DBF" when address_in = 16#04A5# else
		x"2DAE" when address_in = 16#04A6# else
		x"2F2C" when address_in = 16#04A7# else
		x"2F3D" when address_in = 16#04A8# else
		x"2FF3" when address_in = 16#04A9# else
		x"2FE2" when address_in = 16#04AA# else
		x"5AE0" when address_in = 16#04AB# else
		x"4FFF" when address_in = 16#04AC# else
		x"95C8" when address_in = 16#04AD# else
		x"2D80" when address_in = 16#04AE# else
		x"9631" when address_in = 16#04AF# else
		x"95C8" when address_in = 16#04B0# else
		x"2D90" when address_in = 16#04B1# else
		x"938D" when address_in = 16#04B2# else
		x"939D" when address_in = 16#04B3# else
		x"FFC0" when address_in = 16#04B4# else
		x"C003" when address_in = 16#04B5# else
		x"2FF5" when address_in = 16#04B6# else
		x"2FE4" when address_in = 16#04B7# else
		x"C002" when address_in = 16#04B8# else
		x"2FFD" when address_in = 16#04B9# else
		x"2FEC" when address_in = 16#04BA# else
		x"7FEE" when address_in = 16#04BB# else
		x"0FE0" when address_in = 16#04BC# else
		x"1FF1" when address_in = 16#04BD# else
		x"8380" when address_in = 16#04BE# else
		x"8391" when address_in = 16#04BF# else
		x"9621" when address_in = 16#04C0# else
		x"5F2E" when address_in = 16#04C1# else
		x"4F3F" when address_in = 16#04C2# else
		x"5F4F" when address_in = 16#04C3# else
		x"4F5F" when address_in = 16#04C4# else
		x"3FCF" when address_in = 16#04C5# else
		x"05D1" when address_in = 16#04C6# else
		x"F309" when address_in = 16#04C7# else
		x"F304" when address_in = 16#04C8# else
		x"E021" when address_in = 16#04C9# else
		x"BB2B" when address_in = 16#04CA# else
		x"B184" when address_in = 16#04CB# else
		x"2799" when address_in = 16#04CC# else
		x"718E" when address_in = 16#04CD# else
		x"7090" when address_in = 16#04CE# else
		x"9595" when address_in = 16#04CF# else
		x"9587" when address_in = 16#04D0# else
		x"9595" when address_in = 16#04D1# else
		x"9587" when address_in = 16#04D2# else
		x"2F42" when address_in = 16#04D3# else
		x"2F68" when address_in = 16#04D4# else
		x"2F91" when address_in = 16#04D5# else
		x"2F80" when address_in = 16#04D6# else
		x"940E" when address_in = 16#04D7# else
		x"1384" when address_in = 16#04D8# else
		x"E040" when address_in = 16#04D9# else
		x"E050" when address_in = 16#04DA# else
		x"E068" when address_in = 16#04DB# else
		x"E070" when address_in = 16#04DC# else
		x"2F91" when address_in = 16#04DD# else
		x"2F80" when address_in = 16#04DE# else
		x"940E" when address_in = 16#04DF# else
		x"1080" when address_in = 16#04E0# else
		x"E082" when address_in = 16#04E1# else
		x"BB8B" when address_in = 16#04E2# else
		x"E041" when address_in = 16#04E3# else
		x"E050" when address_in = 16#04E4# else
		x"E068" when address_in = 16#04E5# else
		x"E070" when address_in = 16#04E6# else
		x"2F91" when address_in = 16#04E7# else
		x"2F80" when address_in = 16#04E8# else
		x"940E" when address_in = 16#04E9# else
		x"1080" when address_in = 16#04EA# else
		x"2E88" when address_in = 16#04EB# else
		x"2E99" when address_in = 16#04EC# else
		x"E083" when address_in = 16#04ED# else
		x"BB8B" when address_in = 16#04EE# else
		x"E0C0" when address_in = 16#04EF# else
		x"E0D0" when address_in = 16#04F0# else
		x"2DBD" when address_in = 16#04F1# else
		x"2DAC" when address_in = 16#04F2# else
		x"93CD" when address_in = 16#04F3# else
		x"93DC" when address_in = 16#04F4# else
		x"2CAE" when address_in = 16#04F5# else
		x"2CBF" when address_in = 16#04F6# else
		x"2CE1" when address_in = 16#04F7# else
		x"E031" when address_in = 16#04F8# else
		x"2EF3" when address_in = 16#04F9# else
		x"FFC0" when address_in = 16#04FA# else
		x"C003" when address_in = 16#04FB# else
		x"2DFF" when address_in = 16#04FC# else
		x"2DEE" when address_in = 16#04FD# else
		x"C002" when address_in = 16#04FE# else
		x"2FFD" when address_in = 16#04FF# else
		x"2FEC" when address_in = 16#0500# else
		x"7FEE" when address_in = 16#0501# else
		x"0FE0" when address_in = 16#0502# else
		x"1FF1" when address_in = 16#0503# else
		x"9001" when address_in = 16#0504# else
		x"81F0" when address_in = 16#0505# else
		x"2DE0" when address_in = 16#0506# else
		x"2C08" when address_in = 16#0507# else
		x"C002" when address_in = 16#0508# else
		x"0FEE" when address_in = 16#0509# else
		x"1FFF" when address_in = 16#050A# else
		x"940A" when address_in = 16#050B# else
		x"F7E2" when address_in = 16#050C# else
		x"2DBB" when address_in = 16#050D# else
		x"2DAA" when address_in = 16#050E# else
		x"918D" when address_in = 16#050F# else
		x"919D" when address_in = 16#0510# else
		x"2EAA" when address_in = 16#0511# else
		x"2EBB" when address_in = 16#0512# else
		x"1B8E" when address_in = 16#0513# else
		x"0B9F" when address_in = 16#0514# else
		x"940E" when address_in = 16#0515# else
		x"0452" when address_in = 16#0516# else
		x"2DFD" when address_in = 16#0517# else
		x"2DEC" when address_in = 16#0518# else
		x"8120" when address_in = 16#0519# else
		x"8131" when address_in = 16#051A# else
		x"0F28" when address_in = 16#051B# else
		x"1F39" when address_in = 16#051C# else
		x"8320" when address_in = 16#051D# else
		x"8331" when address_in = 16#051E# else
		x"9621" when address_in = 16#051F# else
		x"9408" when address_in = 16#0520# else
		x"1CE1" when address_in = 16#0521# else
		x"1CF1" when address_in = 16#0522# else
		x"3FCF" when address_in = 16#0523# else
		x"05D1" when address_in = 16#0524# else
		x"F2A1" when address_in = 16#0525# else
		x"F29C" when address_in = 16#0526# else
		x"E084" when address_in = 16#0527# else
		x"BB8B" when address_in = 16#0528# else
		x"8180" when address_in = 16#0529# else
		x"BB8B" when address_in = 16#052A# else
		x"8180" when address_in = 16#052B# else
		x"8191" when address_in = 16#052C# else
		x"2F89" when address_in = 16#052D# else
		x"2799" when address_in = 16#052E# else
		x"BB8B" when address_in = 16#052F# else
		x"E085" when address_in = 16#0530# else
		x"BB8B" when address_in = 16#0531# else
		x"CFFF" when address_in = 16#0532# else
		x"93CF" when address_in = 16#0533# else
		x"93DF" when address_in = 16#0534# else
		x"2FF9" when address_in = 16#0535# else
		x"2FE8" when address_in = 16#0536# else
		x"81A2" when address_in = 16#0537# else
		x"81B3" when address_in = 16#0538# else
		x"8184" when address_in = 16#0539# else
		x"8195" when address_in = 16#053A# else
		x"2FDB" when address_in = 16#053B# else
		x"2FCA" when address_in = 16#053C# else
		x"838C" when address_in = 16#053D# else
		x"839D" when address_in = 16#053E# else
		x"8004" when address_in = 16#053F# else
		x"81F5" when address_in = 16#0540# else
		x"2DE0" when address_in = 16#0541# else
		x"83A2" when address_in = 16#0542# else
		x"83B3" when address_in = 16#0543# else
		x"91DF" when address_in = 16#0544# else
		x"91CF" when address_in = 16#0545# else
		x"9508" when address_in = 16#0546# else
		x"EF8F" when address_in = 16#0547# else
		x"BB8B" when address_in = 16#0548# else
		x"B38B" when address_in = 16#0549# else
		x"9580" when address_in = 16#054A# else
		x"CFFC" when address_in = 16#054B# else
		x"93CF" when address_in = 16#054C# else
		x"93DF" when address_in = 16#054D# else
		x"2FF9" when address_in = 16#054E# else
		x"2FE8" when address_in = 16#054F# else
		x"91A0" when address_in = 16#0550# else
		x"0162" when address_in = 16#0551# else
		x"91B0" when address_in = 16#0552# else
		x"0163" when address_in = 16#0553# else
		x"2FDB" when address_in = 16#0554# else
		x"2FCA" when address_in = 16#0555# else
		x"818C" when address_in = 16#0556# else
		x"819D" when address_in = 16#0557# else
		x"83EC" when address_in = 16#0558# else
		x"83FD" when address_in = 16#0559# else
		x"83A2" when address_in = 16#055A# else
		x"83B3" when address_in = 16#055B# else
		x"8384" when address_in = 16#055C# else
		x"8395" when address_in = 16#055D# else
		x"2FD9" when address_in = 16#055E# else
		x"2FC8" when address_in = 16#055F# else
		x"83EA" when address_in = 16#0560# else
		x"83FB" when address_in = 16#0561# else
		x"91DF" when address_in = 16#0562# else
		x"91CF" when address_in = 16#0563# else
		x"9508" when address_in = 16#0564# else
		x"92CF" when address_in = 16#0565# else
		x"92DF" when address_in = 16#0566# else
		x"92EF" when address_in = 16#0567# else
		x"92FF" when address_in = 16#0568# else
		x"930F" when address_in = 16#0569# else
		x"931F" when address_in = 16#056A# else
		x"93CF" when address_in = 16#056B# else
		x"93DF" when address_in = 16#056C# else
		x"2F16" when address_in = 16#056D# else
		x"9700" when address_in = 16#056E# else
		x"F409" when address_in = 16#056F# else
		x"C095" when address_in = 16#0570# else
		x"E059" when address_in = 16#0571# else
		x"2EC5" when address_in = 16#0572# else
		x"2CD1" when address_in = 16#0573# else
		x"0EC8" when address_in = 16#0574# else
		x"1ED9" when address_in = 16#0575# else
		x"E043" when address_in = 16#0576# else
		x"94D6" when address_in = 16#0577# else
		x"94C7" when address_in = 16#0578# else
		x"954A" when address_in = 16#0579# else
		x"F7E1" when address_in = 16#057A# else
		x"B70F" when address_in = 16#057B# else
		x"94F8" when address_in = 16#057C# else
		x"91E0" when address_in = 16#057D# else
		x"0162" when address_in = 16#057E# else
		x"91F0" when address_in = 16#057F# else
		x"0163" when address_in = 16#0580# else
		x"80E4" when address_in = 16#0581# else
		x"80F5" when address_in = 16#0582# else
		x"16EE" when address_in = 16#0583# else
		x"06FF" when address_in = 16#0584# else
		x"F181" when address_in = 16#0585# else
		x"2DBF" when address_in = 16#0586# else
		x"2DAE" when address_in = 16#0587# else
		x"91CD" when address_in = 16#0588# else
		x"91DC" when address_in = 16#0589# else
		x"E033" when address_in = 16#058A# else
		x"0FCC" when address_in = 16#058B# else
		x"1FDD" when address_in = 16#058C# else
		x"953A" when address_in = 16#058D# else
		x"F7E1" when address_in = 16#058E# else
		x"0DCE" when address_in = 16#058F# else
		x"1DDF" when address_in = 16#0590# else
		x"8188" when address_in = 16#0591# else
		x"8199" when address_in = 16#0592# else
		x"2399" when address_in = 16#0593# else
		x"F07C" when address_in = 16#0594# else
		x"2F8C" when address_in = 16#0595# else
		x"2F9D" when address_in = 16#0596# else
		x"940E" when address_in = 16#0597# else
		x"0533" when address_in = 16#0598# else
		x"2DFF" when address_in = 16#0599# else
		x"2DEE" when address_in = 16#059A# else
		x"8180" when address_in = 16#059B# else
		x"8191" when address_in = 16#059C# else
		x"8128" when address_in = 16#059D# else
		x"8139" when address_in = 16#059E# else
		x"0F82" when address_in = 16#059F# else
		x"1F93" when address_in = 16#05A0# else
		x"8380" when address_in = 16#05A1# else
		x"8391" when address_in = 16#05A2# else
		x"CFE2" when address_in = 16#05A3# else
		x"2DBF" when address_in = 16#05A4# else
		x"2DAE" when address_in = 16#05A5# else
		x"918D" when address_in = 16#05A6# else
		x"919C" when address_in = 16#05A7# else
		x"158C" when address_in = 16#05A8# else
		x"059D" when address_in = 16#05A9# else
		x"F458" when address_in = 16#05AA# else
		x"2DFF" when address_in = 16#05AB# else
		x"2DEE" when address_in = 16#05AC# else
		x"80E4" when address_in = 16#05AD# else
		x"80F5" when address_in = 16#05AE# else
		x"9180" when address_in = 16#05AF# else
		x"0162" when address_in = 16#05B0# else
		x"9190" when address_in = 16#05B1# else
		x"0163" when address_in = 16#05B2# else
		x"16E8" when address_in = 16#05B3# else
		x"06F9" when address_in = 16#05B4# else
		x"F681" when address_in = 16#05B5# else
		x"9180" when address_in = 16#05B6# else
		x"0162" when address_in = 16#05B7# else
		x"9190" when address_in = 16#05B8# else
		x"0163" when address_in = 16#05B9# else
		x"16E8" when address_in = 16#05BA# else
		x"06F9" when address_in = 16#05BB# else
		x"F421" when address_in = 16#05BC# else
		x"BF0F" when address_in = 16#05BD# else
		x"E080" when address_in = 16#05BE# else
		x"E090" when address_in = 16#05BF# else
		x"C045" when address_in = 16#05C0# else
		x"2DBF" when address_in = 16#05C1# else
		x"2DAE" when address_in = 16#05C2# else
		x"918D" when address_in = 16#05C3# else
		x"919C" when address_in = 16#05C4# else
		x"9711" when address_in = 16#05C5# else
		x"16C8" when address_in = 16#05C6# else
		x"06D9" when address_in = 16#05C7# else
		x"F498" when address_in = 16#05C8# else
		x"2DFD" when address_in = 16#05C9# else
		x"2DEC" when address_in = 16#05CA# else
		x"E023" when address_in = 16#05CB# else
		x"0FEE" when address_in = 16#05CC# else
		x"1FFF" when address_in = 16#05CD# else
		x"952A" when address_in = 16#05CE# else
		x"F7E1" when address_in = 16#05CF# else
		x"0DEE" when address_in = 16#05D0# else
		x"1DFF" when address_in = 16#05D1# else
		x"198C" when address_in = 16#05D2# else
		x"099D" when address_in = 16#05D3# else
		x"8380" when address_in = 16#05D4# else
		x"8391" when address_in = 16#05D5# else
		x"92CD" when address_in = 16#05D6# else
		x"92DC" when address_in = 16#05D7# else
		x"2F8E" when address_in = 16#05D8# else
		x"2F9F" when address_in = 16#05D9# else
		x"940E" when address_in = 16#05DA# else
		x"054C" when address_in = 16#05DB# else
		x"2D9F" when address_in = 16#05DC# else
		x"2D8E" when address_in = 16#05DD# else
		x"940E" when address_in = 16#05DE# else
		x"0533" when address_in = 16#05DF# else
		x"2DFF" when address_in = 16#05E0# else
		x"2DEE" when address_in = 16#05E1# else
		x"8180" when address_in = 16#05E2# else
		x"8191" when address_in = 16#05E3# else
		x"6890" when address_in = 16#05E4# else
		x"8380" when address_in = 16#05E5# else
		x"8391" when address_in = 16#05E6# else
		x"7017" when address_in = 16#05E7# else
		x"2F81" when address_in = 16#05E8# else
		x"6088" when address_in = 16#05E9# else
		x"2F48" when address_in = 16#05EA# else
		x"E068" when address_in = 16#05EB# else
		x"E070" when address_in = 16#05EC# else
		x"2D9F" when address_in = 16#05ED# else
		x"2D8E" when address_in = 16#05EE# else
		x"940E" when address_in = 16#05EF# else
		x"0797" when address_in = 16#05F0# else
		x"E083" when address_in = 16#05F1# else
		x"0CCC" when address_in = 16#05F2# else
		x"1CDD" when address_in = 16#05F3# else
		x"958A" when address_in = 16#05F4# else
		x"F7E1" when address_in = 16#05F5# else
		x"EF88" when address_in = 16#05F6# else
		x"EF9F" when address_in = 16#05F7# else
		x"0EC8" when address_in = 16#05F8# else
		x"1ED9" when address_in = 16#05F9# else
		x"2F41" when address_in = 16#05FA# else
		x"2D7D" when address_in = 16#05FB# else
		x"2D6C" when address_in = 16#05FC# else
		x"2D9F" when address_in = 16#05FD# else
		x"2D8E" when address_in = 16#05FE# else
		x"9608" when address_in = 16#05FF# else
		x"940E" when address_in = 16#0600# else
		x"0797" when address_in = 16#0601# else
		x"BF0F" when address_in = 16#0602# else
		x"2D9F" when address_in = 16#0603# else
		x"2D8E" when address_in = 16#0604# else
		x"9602" when address_in = 16#0605# else
		x"91DF" when address_in = 16#0606# else
		x"91CF" when address_in = 16#0607# else
		x"911F" when address_in = 16#0608# else
		x"910F" when address_in = 16#0609# else
		x"90FF" when address_in = 16#060A# else
		x"90EF" when address_in = 16#060B# else
		x"90DF" when address_in = 16#060C# else
		x"90CF" when address_in = 16#060D# else
		x"9508" when address_in = 16#060E# else
		x"92EF" when address_in = 16#060F# else
		x"92FF" when address_in = 16#0610# else
		x"931F" when address_in = 16#0611# else
		x"93CF" when address_in = 16#0612# else
		x"93DF" when address_in = 16#0613# else
		x"2EE8" when address_in = 16#0614# else
		x"2EF9" when address_in = 16#0615# else
		x"9700" when address_in = 16#0616# else
		x"F409" when address_in = 16#0617# else
		x"C073" when address_in = 16#0618# else
		x"2FD9" when address_in = 16#0619# else
		x"2FC8" when address_in = 16#061A# else
		x"9722" when address_in = 16#061B# else
		x"E021" when address_in = 16#061C# else
		x"36C8" when address_in = 16#061D# else
		x"07D2" when address_in = 16#061E# else
		x"F408" when address_in = 16#061F# else
		x"C06B" when address_in = 16#0620# else
		x"9180" when address_in = 16#0621# else
		x"0164" when address_in = 16#0622# else
		x"9190" when address_in = 16#0623# else
		x"0165" when address_in = 16#0624# else
		x"E0A3" when address_in = 16#0625# else
		x"0F88" when address_in = 16#0626# else
		x"1F99" when address_in = 16#0627# else
		x"95AA" when address_in = 16#0628# else
		x"F7E1" when address_in = 16#0629# else
		x"5988" when address_in = 16#062A# else
		x"4F9E" when address_in = 16#062B# else
		x"17C8" when address_in = 16#062C# else
		x"07D9" when address_in = 16#062D# else
		x"F008" when address_in = 16#062E# else
		x"C05C" when address_in = 16#062F# else
		x"B71F" when address_in = 16#0630# else
		x"94F8" when address_in = 16#0631# else
		x"B187" when address_in = 16#0632# else
		x"2799" when address_in = 16#0633# else
		x"2F98" when address_in = 16#0634# else
		x"2788" when address_in = 16#0635# else
		x"B128" when address_in = 16#0636# else
		x"2733" when address_in = 16#0637# else
		x"2B82" when address_in = 16#0638# else
		x"2B93" when address_in = 16#0639# else
		x"2F2C" when address_in = 16#063A# else
		x"2F3D" when address_in = 16#063B# else
		x"1B28" when address_in = 16#063C# else
		x"0B39" when address_in = 16#063D# else
		x"2FB3" when address_in = 16#063E# else
		x"2FA2" when address_in = 16#063F# else
		x"95B6" when address_in = 16#0640# else
		x"95A7" when address_in = 16#0641# else
		x"2FF3" when address_in = 16#0642# else
		x"2FE2" when address_in = 16#0643# else
		x"E074" when address_in = 16#0644# else
		x"95F6" when address_in = 16#0645# else
		x"95E7" when address_in = 16#0646# else
		x"957A" when address_in = 16#0647# else
		x"F7E1" when address_in = 16#0648# else
		x"5AE0" when address_in = 16#0649# else
		x"4FFF" when address_in = 16#064A# else
		x"8140" when address_in = 16#064B# else
		x"2F84" when address_in = 16#064C# else
		x"2799" when address_in = 16#064D# else
		x"70A4" when address_in = 16#064E# else
		x"70B0" when address_in = 16#064F# else
		x"2E0A" when address_in = 16#0650# else
		x"C002" when address_in = 16#0651# else
		x"9595" when address_in = 16#0652# else
		x"9587" when address_in = 16#0653# else
		x"940A" when address_in = 16#0654# else
		x"F7E2" when address_in = 16#0655# else
		x"2F48" when address_in = 16#0656# else
		x"704F" when address_in = 16#0657# else
		x"2F24" when address_in = 16#0658# else
		x"2733" when address_in = 16#0659# else
		x"2F93" when address_in = 16#065A# else
		x"2F82" when address_in = 16#065B# else
		x"7088" when address_in = 16#065C# else
		x"7090" when address_in = 16#065D# else
		x"5F87" when address_in = 16#065E# else
		x"4F9F" when address_in = 16#065F# else
		x"F411" when address_in = 16#0660# else
		x"BF1F" when address_in = 16#0661# else
		x"C008" when address_in = 16#0662# else
		x"7027" when address_in = 16#0663# else
		x"7030" when address_in = 16#0664# else
		x"2F86" when address_in = 16#0665# else
		x"2799" when address_in = 16#0666# else
		x"1728" when address_in = 16#0667# else
		x"0739" when address_in = 16#0668# else
		x"F021" when address_in = 16#0669# else
		x"BF1F" when address_in = 16#066A# else
		x"940E" when address_in = 16#066B# else
		x"0547" when address_in = 16#066C# else
		x"C01E" when address_in = 16#066D# else
		x"B71F" when address_in = 16#066E# else
		x"94F8" when address_in = 16#066F# else
		x"8188" when address_in = 16#0670# else
		x"8199" when address_in = 16#0671# else
		x"779F" when address_in = 16#0672# else
		x"8388" when address_in = 16#0673# else
		x"8399" when address_in = 16#0674# else
		x"8120" when address_in = 16#0675# else
		x"E08F" when address_in = 16#0676# else
		x"E090" when address_in = 16#0677# else
		x"C002" when address_in = 16#0678# else
		x"0F88" when address_in = 16#0679# else
		x"1F99" when address_in = 16#067A# else
		x"95AA" when address_in = 16#067B# else
		x"F7E2" when address_in = 16#067C# else
		x"2B28" when address_in = 16#067D# else
		x"8320" when address_in = 16#067E# else
		x"7047" when address_in = 16#067F# else
		x"E02F" when address_in = 16#0680# else
		x"2F62" when address_in = 16#0681# else
		x"2D9F" when address_in = 16#0682# else
		x"2D8E" when address_in = 16#0683# else
		x"9606" when address_in = 16#0684# else
		x"940E" when address_in = 16#0685# else
		x"07F2" when address_in = 16#0686# else
		x"2F8C" when address_in = 16#0687# else
		x"2F9D" when address_in = 16#0688# else
		x"940E" when address_in = 16#0689# else
		x"054C" when address_in = 16#068A# else
		x"BF1F" when address_in = 16#068B# else
		x"91DF" when address_in = 16#068C# else
		x"91CF" when address_in = 16#068D# else
		x"911F" when address_in = 16#068E# else
		x"90FF" when address_in = 16#068F# else
		x"90EF" when address_in = 16#0690# else
		x"9508" when address_in = 16#0691# else
		x"928F" when address_in = 16#0692# else
		x"929F" when address_in = 16#0693# else
		x"92AF" when address_in = 16#0694# else
		x"92BF" when address_in = 16#0695# else
		x"92CF" when address_in = 16#0696# else
		x"92DF" when address_in = 16#0697# else
		x"92EF" when address_in = 16#0698# else
		x"92FF" when address_in = 16#0699# else
		x"930F" when address_in = 16#069A# else
		x"931F" when address_in = 16#069B# else
		x"93CF" when address_in = 16#069C# else
		x"93DF" when address_in = 16#069D# else
		x"2EA8" when address_in = 16#069E# else
		x"2EB9" when address_in = 16#069F# else
		x"2E86" when address_in = 16#06A0# else
		x"2E94" when address_in = 16#06A1# else
		x"2F48" when address_in = 16#06A2# else
		x"2F59" when address_in = 16#06A3# else
		x"5042" when address_in = 16#06A4# else
		x"4050" when address_in = 16#06A5# else
		x"2B89" when address_in = 16#06A6# else
		x"F409" when address_in = 16#06A7# else
		x"C06C" when address_in = 16#06A8# else
		x"B70F" when address_in = 16#06A9# else
		x"94F8" when address_in = 16#06AA# else
		x"B187" when address_in = 16#06AB# else
		x"2799" when address_in = 16#06AC# else
		x"2F98" when address_in = 16#06AD# else
		x"2788" when address_in = 16#06AE# else
		x"B128" when address_in = 16#06AF# else
		x"2733" when address_in = 16#06B0# else
		x"2B82" when address_in = 16#06B1# else
		x"2B93" when address_in = 16#06B2# else
		x"1B48" when address_in = 16#06B3# else
		x"0B59" when address_in = 16#06B4# else
		x"2EE4" when address_in = 16#06B5# else
		x"2EF5" when address_in = 16#06B6# else
		x"94F6" when address_in = 16#06B7# else
		x"94E7" when address_in = 16#06B8# else
		x"2EC4" when address_in = 16#06B9# else
		x"2ED5" when address_in = 16#06BA# else
		x"E0B4" when address_in = 16#06BB# else
		x"94D6" when address_in = 16#06BC# else
		x"94C7" when address_in = 16#06BD# else
		x"95BA" when address_in = 16#06BE# else
		x"F7E1" when address_in = 16#06BF# else
		x"E680" when address_in = 16#06C0# else
		x"E090" when address_in = 16#06C1# else
		x"0EC8" when address_in = 16#06C2# else
		x"1ED9" when address_in = 16#06C3# else
		x"2DFD" when address_in = 16#06C4# else
		x"2DEC" when address_in = 16#06C5# else
		x"8110" when address_in = 16#06C6# else
		x"2F81" when address_in = 16#06C7# else
		x"2799" when address_in = 16#06C8# else
		x"E0F4" when address_in = 16#06C9# else
		x"22EF" when address_in = 16#06CA# else
		x"24FF" when address_in = 16#06CB# else
		x"2C0E" when address_in = 16#06CC# else
		x"C002" when address_in = 16#06CD# else
		x"9595" when address_in = 16#06CE# else
		x"9587" when address_in = 16#06CF# else
		x"940A" when address_in = 16#06D0# else
		x"F7E2" when address_in = 16#06D1# else
		x"2F18" when address_in = 16#06D2# else
		x"701F" when address_in = 16#06D3# else
		x"2FC1" when address_in = 16#06D4# else
		x"27DD" when address_in = 16#06D5# else
		x"2F8C" when address_in = 16#06D6# else
		x"2F9D" when address_in = 16#06D7# else
		x"7088" when address_in = 16#06D8# else
		x"7090" when address_in = 16#06D9# else
		x"5F87" when address_in = 16#06DA# else
		x"4F9F" when address_in = 16#06DB# else
		x"F419" when address_in = 16#06DC# else
		x"BF0F" when address_in = 16#06DD# else
		x"940E" when address_in = 16#06DE# else
		x"0547" when address_in = 16#06DF# else
		x"2F2C" when address_in = 16#06E0# else
		x"2F3D" when address_in = 16#06E1# else
		x"7027" when address_in = 16#06E2# else
		x"7030" when address_in = 16#06E3# else
		x"2D88" when address_in = 16#06E4# else
		x"2799" when address_in = 16#06E5# else
		x"1728" when address_in = 16#06E6# else
		x"0739" when address_in = 16#06E7# else
		x"F549" when address_in = 16#06E8# else
		x"2D49" when address_in = 16#06E9# else
		x"2755" when address_in = 16#06EA# else
		x"1742" when address_in = 16#06EB# else
		x"0753" when address_in = 16#06EC# else
		x"F151" when address_in = 16#06ED# else
		x"2DFD" when address_in = 16#06EE# else
		x"2DEC" when address_in = 16#06EF# else
		x"8180" when address_in = 16#06F0# else
		x"E02F" when address_in = 16#06F1# else
		x"E030" when address_in = 16#06F2# else
		x"2C0E" when address_in = 16#06F3# else
		x"C002" when address_in = 16#06F4# else
		x"0F22" when address_in = 16#06F5# else
		x"1F33" when address_in = 16#06F6# else
		x"940A" when address_in = 16#06F7# else
		x"F7E2" when address_in = 16#06F8# else
		x"2F92" when address_in = 16#06F9# else
		x"9590" when address_in = 16#06FA# else
		x"2389" when address_in = 16#06FB# else
		x"7047" when address_in = 16#06FC# else
		x"7050" when address_in = 16#06FD# else
		x"6048" when address_in = 16#06FE# else
		x"C002" when address_in = 16#06FF# else
		x"0F44" when address_in = 16#0700# else
		x"1F55" when address_in = 16#0701# else
		x"94EA" when address_in = 16#0702# else
		x"F7E2" when address_in = 16#0703# else
		x"2B84" when address_in = 16#0704# else
		x"8380" when address_in = 16#0705# else
		x"E0F7" when address_in = 16#0706# else
		x"229F" when address_in = 16#0707# else
		x"231F" when address_in = 16#0708# else
		x"2D29" when address_in = 16#0709# else
		x"2F41" when address_in = 16#070A# else
		x"E06F" when address_in = 16#070B# else
		x"2D9B" when address_in = 16#070C# else
		x"2D8A" when address_in = 16#070D# else
		x"9606" when address_in = 16#070E# else
		x"940E" when address_in = 16#070F# else
		x"07F2" when address_in = 16#0710# else
		x"C006" when address_in = 16#0711# else
		x"BF0F" when address_in = 16#0712# else
		x"940E" when address_in = 16#0713# else
		x"0547" when address_in = 16#0714# else
		x"EF8F" when address_in = 16#0715# else
		x"EF9F" when address_in = 16#0716# else
		x"C003" when address_in = 16#0717# else
		x"BF0F" when address_in = 16#0718# else
		x"E080" when address_in = 16#0719# else
		x"E090" when address_in = 16#071A# else
		x"91DF" when address_in = 16#071B# else
		x"91CF" when address_in = 16#071C# else
		x"911F" when address_in = 16#071D# else
		x"910F" when address_in = 16#071E# else
		x"90FF" when address_in = 16#071F# else
		x"90EF" when address_in = 16#0720# else
		x"90DF" when address_in = 16#0721# else
		x"90CF" when address_in = 16#0722# else
		x"90BF" when address_in = 16#0723# else
		x"90AF" when address_in = 16#0724# else
		x"909F" when address_in = 16#0725# else
		x"908F" when address_in = 16#0726# else
		x"9508" when address_in = 16#0727# else
		x"92EF" when address_in = 16#0728# else
		x"92FF" when address_in = 16#0729# else
		x"930F" when address_in = 16#072A# else
		x"931F" when address_in = 16#072B# else
		x"E608" when address_in = 16#072C# else
		x"E011" when address_in = 16#072D# else
		x"2CE1" when address_in = 16#072E# else
		x"E038" when address_in = 16#072F# else
		x"2EF3" when address_in = 16#0730# else
		x"0EE0" when address_in = 16#0731# else
		x"1EF1" when address_in = 16#0732# else
		x"9310" when address_in = 16#0733# else
		x"0161" when address_in = 16#0734# else
		x"9300" when address_in = 16#0735# else
		x"0160" when address_in = 16#0736# else
		x"EF4F" when address_in = 16#0737# else
		x"E050" when address_in = 16#0738# else
		x"9350" when address_in = 16#0739# else
		x"0165" when address_in = 16#073A# else
		x"9340" when address_in = 16#073B# else
		x"0164" when address_in = 16#073C# else
		x"2F31" when address_in = 16#073D# else
		x"2F20" when address_in = 16#073E# else
		x"5028" when address_in = 16#073F# else
		x"4F38" when address_in = 16#0740# else
		x"9330" when address_in = 16#0741# else
		x"0163" when address_in = 16#0742# else
		x"9320" when address_in = 16#0743# else
		x"0162" when address_in = 16#0744# else
		x"E080" when address_in = 16#0745# else
		x"E890" when address_in = 16#0746# else
		x"9390" when address_in = 16#0747# else
		x"0961" when address_in = 16#0748# else
		x"9380" when address_in = 16#0749# else
		x"0960" when address_in = 16#074A# else
		x"9330" when address_in = 16#074B# else
		x"0963" when address_in = 16#074C# else
		x"9320" when address_in = 16#074D# else
		x"0962" when address_in = 16#074E# else
		x"9330" when address_in = 16#074F# else
		x"0965" when address_in = 16#0750# else
		x"9320" when address_in = 16#0751# else
		x"0964" when address_in = 16#0752# else
		x"9350" when address_in = 16#0753# else
		x"0169" when address_in = 16#0754# else
		x"9340" when address_in = 16#0755# else
		x"0168" when address_in = 16#0756# else
		x"2F91" when address_in = 16#0757# else
		x"2F80" when address_in = 16#0758# else
		x"940E" when address_in = 16#0759# else
		x"054C" when address_in = 16#075A# else
		x"940E" when address_in = 16#075B# else
		x"078D" when address_in = 16#075C# else
		x"9180" when address_in = 16#075D# else
		x"0164" when address_in = 16#075E# else
		x"9190" when address_in = 16#075F# else
		x"0165" when address_in = 16#0760# else
		x"E023" when address_in = 16#0761# else
		x"0F88" when address_in = 16#0762# else
		x"1F99" when address_in = 16#0763# else
		x"952A" when address_in = 16#0764# else
		x"F7E1" when address_in = 16#0765# else
		x"E04F" when address_in = 16#0766# else
		x"2F68" when address_in = 16#0767# else
		x"2F79" when address_in = 16#0768# else
		x"9180" when address_in = 16#0769# else
		x"0160" when address_in = 16#076A# else
		x"9190" when address_in = 16#076B# else
		x"0161" when address_in = 16#076C# else
		x"940E" when address_in = 16#076D# else
		x"0797" when address_in = 16#076E# else
		x"B184" when address_in = 16#076F# else
		x"718F" when address_in = 16#0770# else
		x"B984" when address_in = 16#0771# else
		x"B184" when address_in = 16#0772# else
		x"6680" when address_in = 16#0773# else
		x"B984" when address_in = 16#0774# else
		x"9821" when address_in = 16#0775# else
		x"B908" when address_in = 16#0776# else
		x"2F81" when address_in = 16#0777# else
		x"2799" when address_in = 16#0778# else
		x"B987" when address_in = 16#0779# else
		x"B8E6" when address_in = 16#077A# else
		x"2D8F" when address_in = 16#077B# else
		x"2799" when address_in = 16#077C# else
		x"B985" when address_in = 16#077D# else
		x"E680" when address_in = 16#077E# else
		x"E090" when address_in = 16#077F# else
		x"BB8D" when address_in = 16#0780# else
		x"2F89" when address_in = 16#0781# else
		x"2799" when address_in = 16#0782# else
		x"BB8E" when address_in = 16#0783# else
		x"BA1C" when address_in = 16#0784# else
		x"E180" when address_in = 16#0785# else
		x"BB8F" when address_in = 16#0786# else
		x"9A20" when address_in = 16#0787# else
		x"911F" when address_in = 16#0788# else
		x"910F" when address_in = 16#0789# else
		x"90FF" when address_in = 16#078A# else
		x"90EF" when address_in = 16#078B# else
		x"9508" when address_in = 16#078C# else
		x"EF8F" when address_in = 16#078D# else
		x"E6E0" when address_in = 16#078E# else
		x"E0F0" when address_in = 16#078F# else
		x"9381" when address_in = 16#0790# else
		x"E091" when address_in = 16#0791# else
		x"35EF" when address_in = 16#0792# else
		x"07F9" when address_in = 16#0793# else
		x"F3D9" when address_in = 16#0794# else
		x"F3D0" when address_in = 16#0795# else
		x"9508" when address_in = 16#0796# else
		x"93CF" when address_in = 16#0797# else
		x"2FF9" when address_in = 16#0798# else
		x"2FE8" when address_in = 16#0799# else
		x"2FC4" when address_in = 16#079A# else
		x"1561" when address_in = 16#079B# else
		x"0571" when address_in = 16#079C# else
		x"F409" when address_in = 16#079D# else
		x"C051" when address_in = 16#079E# else
		x"2F97" when address_in = 16#079F# else
		x"2F86" when address_in = 16#07A0# else
		x"7087" when address_in = 16#07A1# else
		x"7F98" when address_in = 16#07A2# else
		x"2B89" when address_in = 16#07A3# else
		x"F009" when address_in = 16#07A4# else
		x"C04A" when address_in = 16#07A5# else
		x"E043" when address_in = 16#07A6# else
		x"9576" when address_in = 16#07A7# else
		x"9567" when address_in = 16#07A8# else
		x"954A" when address_in = 16#07A9# else
		x"F7E1" when address_in = 16#07AA# else
		x"B187" when address_in = 16#07AB# else
		x"2799" when address_in = 16#07AC# else
		x"2F98" when address_in = 16#07AD# else
		x"2788" when address_in = 16#07AE# else
		x"B128" when address_in = 16#07AF# else
		x"2733" when address_in = 16#07B0# else
		x"2B82" when address_in = 16#07B1# else
		x"2B93" when address_in = 16#07B2# else
		x"1BE8" when address_in = 16#07B3# else
		x"0BF9" when address_in = 16#07B4# else
		x"2FAE" when address_in = 16#07B5# else
		x"2FBF" when address_in = 16#07B6# else
		x"E024" when address_in = 16#07B7# else
		x"95B6" when address_in = 16#07B8# else
		x"95A7" when address_in = 16#07B9# else
		x"952A" when address_in = 16#07BA# else
		x"F7E1" when address_in = 16#07BB# else
		x"2F2E" when address_in = 16#07BC# else
		x"2F3F" when address_in = 16#07BD# else
		x"9536" when address_in = 16#07BE# else
		x"9527" when address_in = 16#07BF# else
		x"2FFB" when address_in = 16#07C0# else
		x"2FEA" when address_in = 16#07C1# else
		x"5AE0" when address_in = 16#07C2# else
		x"4FFF" when address_in = 16#07C3# else
		x"8150" when address_in = 16#07C4# else
		x"7024" when address_in = 16#07C5# else
		x"7030" when address_in = 16#07C6# else
		x"E08F" when address_in = 16#07C7# else
		x"E090" when address_in = 16#07C8# else
		x"2E02" when address_in = 16#07C9# else
		x"C002" when address_in = 16#07CA# else
		x"0F88" when address_in = 16#07CB# else
		x"1F99" when address_in = 16#07CC# else
		x"940A" when address_in = 16#07CD# else
		x"F7E2" when address_in = 16#07CE# else
		x"2F48" when address_in = 16#07CF# else
		x"2F8C" when address_in = 16#07D0# else
		x"2799" when address_in = 16#07D1# else
		x"C002" when address_in = 16#07D2# else
		x"0F88" when address_in = 16#07D3# else
		x"1F99" when address_in = 16#07D4# else
		x"952A" when address_in = 16#07D5# else
		x"F7E2" when address_in = 16#07D6# else
		x"2F98" when address_in = 16#07D7# else
		x"1561" when address_in = 16#07D8# else
		x"0571" when address_in = 16#07D9# else
		x"F091" when address_in = 16#07DA# else
		x"2F84" when address_in = 16#07DB# else
		x"9580" when address_in = 16#07DC# else
		x"2358" when address_in = 16#07DD# else
		x"2B59" when address_in = 16#07DE# else
		x"5061" when address_in = 16#07DF# else
		x"4070" when address_in = 16#07E0# else
		x"9542" when address_in = 16#07E1# else
		x"7F40" when address_in = 16#07E2# else
		x"9592" when address_in = 16#07E3# else
		x"7F90" when address_in = 16#07E4# else
		x"2344" when address_in = 16#07E5# else
		x"F789" when address_in = 16#07E6# else
		x"9351" when address_in = 16#07E7# else
		x"9611" when address_in = 16#07E8# else
		x"8150" when address_in = 16#07E9# else
		x"E04F" when address_in = 16#07EA# else
		x"2F9C" when address_in = 16#07EB# else
		x"CFEB" when address_in = 16#07EC# else
		x"5AA0" when address_in = 16#07ED# else
		x"4FBF" when address_in = 16#07EE# else
		x"935C" when address_in = 16#07EF# else
		x"91CF" when address_in = 16#07F0# else
		x"9508" when address_in = 16#07F1# else
		x"92FF" when address_in = 16#07F2# else
		x"930F" when address_in = 16#07F3# else
		x"931F" when address_in = 16#07F4# else
		x"93CF" when address_in = 16#07F5# else
		x"93DF" when address_in = 16#07F6# else
		x"2EF6" when address_in = 16#07F7# else
		x"2F04" when address_in = 16#07F8# else
		x"2F12" when address_in = 16#07F9# else
		x"E0C0" when address_in = 16#07FA# else
		x"E0D0" when address_in = 16#07FB# else
		x"B127" when address_in = 16#07FC# else
		x"2733" when address_in = 16#07FD# else
		x"2F32" when address_in = 16#07FE# else
		x"2722" when address_in = 16#07FF# else
		x"B148" when address_in = 16#0800# else
		x"2755" when address_in = 16#0801# else
		x"2B24" when address_in = 16#0802# else
		x"2B35" when address_in = 16#0803# else
		x"1B82" when address_in = 16#0804# else
		x"0B93" when address_in = 16#0805# else
		x"2FB9" when address_in = 16#0806# else
		x"2FA8" when address_in = 16#0807# else
		x"E064" when address_in = 16#0808# else
		x"95B6" when address_in = 16#0809# else
		x"95A7" when address_in = 16#080A# else
		x"956A" when address_in = 16#080B# else
		x"F7E1" when address_in = 16#080C# else
		x"2F28" when address_in = 16#080D# else
		x"2F39" when address_in = 16#080E# else
		x"9536" when address_in = 16#080F# else
		x"9527" when address_in = 16#0810# else
		x"2FFB" when address_in = 16#0811# else
		x"2FEA" when address_in = 16#0812# else
		x"5AE0" when address_in = 16#0813# else
		x"4FFF" when address_in = 16#0814# else
		x"8140" when address_in = 16#0815# else
		x"2D8F" when address_in = 16#0816# else
		x"2799" when address_in = 16#0817# else
		x"7024" when address_in = 16#0818# else
		x"7030" when address_in = 16#0819# else
		x"2E02" when address_in = 16#081A# else
		x"C002" when address_in = 16#081B# else
		x"0F88" when address_in = 16#081C# else
		x"1F99" when address_in = 16#081D# else
		x"940A" when address_in = 16#081E# else
		x"F7E2" when address_in = 16#081F# else
		x"2F68" when address_in = 16#0820# else
		x"2F80" when address_in = 16#0821# else
		x"2799" when address_in = 16#0822# else
		x"2E02" when address_in = 16#0823# else
		x"C002" when address_in = 16#0824# else
		x"0F88" when address_in = 16#0825# else
		x"1F99" when address_in = 16#0826# else
		x"940A" when address_in = 16#0827# else
		x"F7E2" when address_in = 16#0828# else
		x"2F58" when address_in = 16#0829# else
		x"2F81" when address_in = 16#082A# else
		x"2799" when address_in = 16#082B# else
		x"2E02" when address_in = 16#082C# else
		x"C002" when address_in = 16#082D# else
		x"0F88" when address_in = 16#082E# else
		x"1F99" when address_in = 16#082F# else
		x"940A" when address_in = 16#0830# else
		x"F7E2" when address_in = 16#0831# else
		x"2F78" when address_in = 16#0832# else
		x"E08F" when address_in = 16#0833# else
		x"E090" when address_in = 16#0834# else
		x"C002" when address_in = 16#0835# else
		x"0F88" when address_in = 16#0836# else
		x"1F99" when address_in = 16#0837# else
		x"952A" when address_in = 16#0838# else
		x"F7E2" when address_in = 16#0839# else
		x"2F98" when address_in = 16#083A# else
		x"2F84" when address_in = 16#083B# else
		x"2386" when address_in = 16#083C# else
		x"1785" when address_in = 16#083D# else
		x"F4B1" when address_in = 16#083E# else
		x"2F89" when address_in = 16#083F# else
		x"9580" when address_in = 16#0840# else
		x"2348" when address_in = 16#0841# else
		x"2B47" when address_in = 16#0842# else
		x"9621" when address_in = 16#0843# else
		x"9562" when address_in = 16#0844# else
		x"7F60" when address_in = 16#0845# else
		x"9552" when address_in = 16#0846# else
		x"7F50" when address_in = 16#0847# else
		x"9572" when address_in = 16#0848# else
		x"7F70" when address_in = 16#0849# else
		x"9592" when address_in = 16#084A# else
		x"7F90" when address_in = 16#084B# else
		x"F771" when address_in = 16#084C# else
		x"9341" when address_in = 16#084D# else
		x"9611" when address_in = 16#084E# else
		x"8140" when address_in = 16#084F# else
		x"2D6F" when address_in = 16#0850# else
		x"2F50" when address_in = 16#0851# else
		x"2F71" when address_in = 16#0852# else
		x"E09F" when address_in = 16#0853# else
		x"CFE6" when address_in = 16#0854# else
		x"5AA0" when address_in = 16#0855# else
		x"4FBF" when address_in = 16#0856# else
		x"934C" when address_in = 16#0857# else
		x"2F8C" when address_in = 16#0858# else
		x"2F9D" when address_in = 16#0859# else
		x"91DF" when address_in = 16#085A# else
		x"91CF" when address_in = 16#085B# else
		x"911F" when address_in = 16#085C# else
		x"910F" when address_in = 16#085D# else
		x"90FF" when address_in = 16#085E# else
		x"9508" when address_in = 16#085F# else
		x"940E" when address_in = 16#0860# else
		x"0B02" when address_in = 16#0861# else
		x"0F99" when address_in = 16#0862# else
		x"0B88" when address_in = 16#0863# else
		x"0F99" when address_in = 16#0864# else
		x"2F98" when address_in = 16#0865# else
		x"1F88" when address_in = 16#0866# else
		x"2F28" when address_in = 16#0867# else
		x"2F39" when address_in = 16#0868# else
		x"9535" when address_in = 16#0869# else
		x"9527" when address_in = 16#086A# else
		x"7081" when address_in = 16#086B# else
		x"7090" when address_in = 16#086C# else
		x"0F82" when address_in = 16#086D# else
		x"1F93" when address_in = 16#086E# else
		x"9508" when address_in = 16#086F# else
		x"922F" when address_in = 16#0870# else
		x"923F" when address_in = 16#0871# else
		x"924F" when address_in = 16#0872# else
		x"925F" when address_in = 16#0873# else
		x"926F" when address_in = 16#0874# else
		x"927F" when address_in = 16#0875# else
		x"928F" when address_in = 16#0876# else
		x"929F" when address_in = 16#0877# else
		x"92AF" when address_in = 16#0878# else
		x"92BF" when address_in = 16#0879# else
		x"92CF" when address_in = 16#087A# else
		x"92DF" when address_in = 16#087B# else
		x"92EF" when address_in = 16#087C# else
		x"92FF" when address_in = 16#087D# else
		x"930F" when address_in = 16#087E# else
		x"931F" when address_in = 16#087F# else
		x"93CF" when address_in = 16#0880# else
		x"93DF" when address_in = 16#0881# else
		x"B7CD" when address_in = 16#0882# else
		x"B7DE" when address_in = 16#0883# else
		x"9768" when address_in = 16#0884# else
		x"B60F" when address_in = 16#0885# else
		x"94F8" when address_in = 16#0886# else
		x"BFDE" when address_in = 16#0887# else
		x"BE0F" when address_in = 16#0888# else
		x"BFCD" when address_in = 16#0889# else
		x"8389" when address_in = 16#088A# else
		x"839A" when address_in = 16#088B# else
		x"836B" when address_in = 16#088C# else
		x"837C" when address_in = 16#088D# else
		x"8B4D" when address_in = 16#088E# else
		x"8B5E" when address_in = 16#088F# else
		x"832D" when address_in = 16#0890# else
		x"833E" when address_in = 16#0891# else
		x"E081" when address_in = 16#0892# else
		x"E090" when address_in = 16#0893# else
		x"2E68" when address_in = 16#0894# else
		x"2E79" when address_in = 16#0895# else
		x"880D" when address_in = 16#0896# else
		x"C002" when address_in = 16#0897# else
		x"0C66" when address_in = 16#0898# else
		x"1C77" when address_in = 16#0899# else
		x"940A" when address_in = 16#089A# else
		x"F7E2" when address_in = 16#089B# else
		x"E021" when address_in = 16#089C# else
		x"1662" when address_in = 16#089D# else
		x"E024" when address_in = 16#089E# else
		x"0672" when address_in = 16#089F# else
		x"F01C" when address_in = 16#08A0# else
		x"EF8F" when address_in = 16#08A1# else
		x"EF9F" when address_in = 16#08A2# else
		x"C1D5" when address_in = 16#08A3# else
		x"E040" when address_in = 16#08A4# else
		x"E050" when address_in = 16#08A5# else
		x"2CB7" when address_in = 16#08A6# else
		x"2CA6" when address_in = 16#08A7# else
		x"9408" when address_in = 16#08A8# else
		x"08A1" when address_in = 16#08A9# else
		x"08B1" when address_in = 16#08AA# else
		x"874B" when address_in = 16#08AB# else
		x"875C" when address_in = 16#08AC# else
		x"8B8D" when address_in = 16#08AD# else
		x"8B9E" when address_in = 16#08AE# else
		x"16A8" when address_in = 16#08AF# else
		x"06B9" when address_in = 16#08B0# else
		x"F40C" when address_in = 16#08B1# else
		x"C058" when address_in = 16#08B2# else
		x"80EB" when address_in = 16#08B3# else
		x"80FC" when address_in = 16#08B4# else
		x"E082" when address_in = 16#08B5# else
		x"E090" when address_in = 16#08B6# else
		x"0EE8" when address_in = 16#08B7# else
		x"1EF9" when address_in = 16#08B8# else
		x"8169" when address_in = 16#08B9# else
		x"817A" when address_in = 16#08BA# else
		x"0F68" when address_in = 16#08BB# else
		x"1F79" when address_in = 16#08BC# else
		x"2CD7" when address_in = 16#08BD# else
		x"2CC6" when address_in = 16#08BE# else
		x"94D5" when address_in = 16#08BF# else
		x"94C7" when address_in = 16#08C0# else
		x"2F95" when address_in = 16#08C1# else
		x"2F84" when address_in = 16#08C2# else
		x"0D8C" when address_in = 16#08C3# else
		x"1D9D" when address_in = 16#08C4# else
		x"16A8" when address_in = 16#08C5# else
		x"06B9" when address_in = 16#08C6# else
		x"F3BC" when address_in = 16#08C7# else
		x"2D9D" when address_in = 16#08C8# else
		x"2D8C" when address_in = 16#08C9# else
		x"9701" when address_in = 16#08CA# else
		x"2348" when address_in = 16#08CB# else
		x"2359" when address_in = 16#08CC# else
		x"0D4C" when address_in = 16#08CD# else
		x"1D5D" when address_in = 16#08CE# else
		x"89ED" when address_in = 16#08CF# else
		x"89FE" when address_in = 16#08D0# else
		x"17E4" when address_in = 16#08D1# else
		x"07F5" when address_in = 16#08D2# else
		x"F53C" when address_in = 16#08D3# else
		x"2FF7" when address_in = 16#08D4# else
		x"2FE6" when address_in = 16#08D5# else
		x"8100" when address_in = 16#08D6# else
		x"8111" when address_in = 16#08D7# else
		x"2F24" when address_in = 16#08D8# else
		x"2F35" when address_in = 16#08D9# else
		x"0F24" when address_in = 16#08DA# else
		x"1F35" when address_in = 16#08DB# else
		x"81A9" when address_in = 16#08DC# else
		x"81BA" when address_in = 16#08DD# else
		x"0FA2" when address_in = 16#08DE# else
		x"1FB3" when address_in = 16#08DF# else
		x"918D" when address_in = 16#08E0# else
		x"919C" when address_in = 16#08E1# else
		x"9711" when address_in = 16#08E2# else
		x"8380" when address_in = 16#08E3# else
		x"8391" when address_in = 16#08E4# else
		x"930D" when address_in = 16#08E5# else
		x"931C" when address_in = 16#08E6# else
		x"2DFF" when address_in = 16#08E7# else
		x"2DEE" when address_in = 16#08E8# else
		x"81A0" when address_in = 16#08E9# else
		x"81B1" when address_in = 16#08EA# else
		x"818B" when address_in = 16#08EB# else
		x"819C" when address_in = 16#08EC# else
		x"0F28" when address_in = 16#08ED# else
		x"1F39" when address_in = 16#08EE# else
		x"2FF3" when address_in = 16#08EF# else
		x"2FE2" when address_in = 16#08F0# else
		x"8180" when address_in = 16#08F1# else
		x"8191" when address_in = 16#08F2# else
		x"2DFF" when address_in = 16#08F3# else
		x"2DEE" when address_in = 16#08F4# else
		x"8380" when address_in = 16#08F5# else
		x"8391" when address_in = 16#08F6# else
		x"2FF3" when address_in = 16#08F7# else
		x"2FE2" when address_in = 16#08F8# else
		x"83A0" when address_in = 16#08F9# else
		x"83B1" when address_in = 16#08FA# else
		x"892D" when address_in = 16#08FB# else
		x"893E" when address_in = 16#08FC# else
		x"5F2F" when address_in = 16#08FD# else
		x"4F3F" when address_in = 16#08FE# else
		x"8B2D" when address_in = 16#08FF# else
		x"8B3E" when address_in = 16#0900# else
		x"5F6E" when address_in = 16#0901# else
		x"4F7F" when address_in = 16#0902# else
		x"E082" when address_in = 16#0903# else
		x"E090" when address_in = 16#0904# else
		x"0EE8" when address_in = 16#0905# else
		x"1EF9" when address_in = 16#0906# else
		x"16A2" when address_in = 16#0907# else
		x"06B3" when address_in = 16#0908# else
		x"F00C" when address_in = 16#0909# else
		x"CFB2" when address_in = 16#090A# else
		x"E0E1" when address_in = 16#090B# else
		x"2ECE" when address_in = 16#090C# else
		x"2CD1" when address_in = 16#090D# else
		x"E0E9" when address_in = 16#090E# else
		x"E0F0" when address_in = 16#090F# else
		x"83EF" when address_in = 16#0910# else
		x"87F8" when address_in = 16#0911# else
		x"14C6" when address_in = 16#0912# else
		x"04D7" when address_in = 16#0913# else
		x"F00C" when address_in = 16#0914# else
		x"C161" when address_in = 16#0915# else
		x"812D" when address_in = 16#0916# else
		x"813E" when address_in = 16#0917# else
		x"2B23" when address_in = 16#0918# else
		x"F1E1" when address_in = 16#0919# else
		x"24AA" when address_in = 16#091A# else
		x"24BB" when address_in = 16#091B# else
		x"86AD" when address_in = 16#091C# else
		x"86BE" when address_in = 16#091D# else
		x"14A6" when address_in = 16#091E# else
		x"04B7" when address_in = 16#091F# else
		x"F5CC" when address_in = 16#0920# else
		x"814B" when address_in = 16#0921# else
		x"815C" when address_in = 16#0922# else
		x"81A9" when address_in = 16#0923# else
		x"81BA" when address_in = 16#0924# else
		x"918D" when address_in = 16#0925# else
		x"919D" when address_in = 16#0926# else
		x"FF97" when address_in = 16#0927# else
		x"C003" when address_in = 16#0928# else
		x"9590" when address_in = 16#0929# else
		x"9581" when address_in = 16#092A# else
		x"4F9F" when address_in = 16#092B# else
		x"2FF5" when address_in = 16#092C# else
		x"2FE4" when address_in = 16#092D# else
		x"9001" when address_in = 16#092E# else
		x"81F0" when address_in = 16#092F# else
		x"2DE0" when address_in = 16#0930# else
		x"8BED" when address_in = 16#0931# else
		x"8BFE" when address_in = 16#0932# else
		x"FFF7" when address_in = 16#0933# else
		x"C005" when address_in = 16#0934# else
		x"95F0" when address_in = 16#0935# else
		x"95E1" when address_in = 16#0936# else
		x"4FFF" when address_in = 16#0937# else
		x"8BED" when address_in = 16#0938# else
		x"8BFE" when address_in = 16#0939# else
		x"5080" when address_in = 16#093A# else
		x"4490" when address_in = 16#093B# else
		x"F42C" when address_in = 16#093C# else
		x"892D" when address_in = 16#093D# else
		x"893E" when address_in = 16#093E# else
		x"5020" when address_in = 16#093F# else
		x"4430" when address_in = 16#0940# else
		x"F05C" when address_in = 16#0941# else
		x"E0E1" when address_in = 16#0942# else
		x"E0F0" when address_in = 16#0943# else
		x"87ED" when address_in = 16#0944# else
		x"87FE" when address_in = 16#0945# else
		x"852B" when address_in = 16#0946# else
		x"853C" when address_in = 16#0947# else
		x"0F2E" when address_in = 16#0948# else
		x"1F3F" when address_in = 16#0949# else
		x"872B" when address_in = 16#094A# else
		x"873C" when address_in = 16#094B# else
		x"C00D" when address_in = 16#094C# else
		x"9408" when address_in = 16#094D# else
		x"1CA1" when address_in = 16#094E# else
		x"1CB1" when address_in = 16#094F# else
		x"5F4E" when address_in = 16#0950# else
		x"4F5F" when address_in = 16#0951# else
		x"14A6" when address_in = 16#0952# else
		x"04B7" when address_in = 16#0953# else
		x"F284" when address_in = 16#0954# else
		x"C004" when address_in = 16#0955# else
		x"E081" when address_in = 16#0956# else
		x"E090" when address_in = 16#0957# else
		x"878D" when address_in = 16#0958# else
		x"879E" when address_in = 16#0959# else
		x"2DFD" when address_in = 16#095A# else
		x"2DEC" when address_in = 16#095B# else
		x"0FEE" when address_in = 16#095C# else
		x"1FFF" when address_in = 16#095D# else
		x"87E9" when address_in = 16#095E# else
		x"87FA" when address_in = 16#095F# else
		x"8A1D" when address_in = 16#0960# else
		x"8A1E" when address_in = 16#0961# else
		x"E020" when address_in = 16#0962# else
		x"E030" when address_in = 16#0963# else
		x"152C" when address_in = 16#0964# else
		x"053D" when address_in = 16#0965# else
		x"F00C" when address_in = 16#0966# else
		x"C107" when address_in = 16#0967# else
		x"8B2B" when address_in = 16#0968# else
		x"8B3C" when address_in = 16#0969# else
		x"898D" when address_in = 16#096A# else
		x"899E" when address_in = 16#096B# else
		x"800F" when address_in = 16#096C# else
		x"C002" when address_in = 16#096D# else
		x"0F88" when address_in = 16#096E# else
		x"1F99" when address_in = 16#096F# else
		x"940A" when address_in = 16#0970# else
		x"F7E2" when address_in = 16#0971# else
		x"0F88" when address_in = 16#0972# else
		x"1F99" when address_in = 16#0973# else
		x"2F68" when address_in = 16#0974# else
		x"2F79" when address_in = 16#0975# else
		x"5A60" when address_in = 16#0976# else
		x"4F7B" when address_in = 16#0977# else
		x"2FF7" when address_in = 16#0978# else
		x"2FE6" when address_in = 16#0979# else
		x"95C8" when address_in = 16#097A# else
		x"2D20" when address_in = 16#097B# else
		x"9631" when address_in = 16#097C# else
		x"95C8" when address_in = 16#097D# else
		x"2D30" when address_in = 16#097E# else
		x"872F" when address_in = 16#097F# else
		x"8B38" when address_in = 16#0980# else
		x"2FF9" when address_in = 16#0981# else
		x"2FE8" when address_in = 16#0982# else
		x"5AE0" when address_in = 16#0983# else
		x"4FFD" when address_in = 16#0984# else
		x"95C8" when address_in = 16#0985# else
		x"2D80" when address_in = 16#0986# else
		x"9631" when address_in = 16#0987# else
		x"95C8" when address_in = 16#0988# else
		x"2D90" when address_in = 16#0989# else
		x"2444" when address_in = 16#098A# else
		x"2455" when address_in = 16#098B# else
		x"1A48" when address_in = 16#098C# else
		x"0A59" when address_in = 16#098D# else
		x"81ED" when address_in = 16#098E# else
		x"81FE" when address_in = 16#098F# else
		x"2BEF" when address_in = 16#0990# else
		x"F011" when address_in = 16#0991# else
		x"2E48" when address_in = 16#0992# else
		x"2E59" when address_in = 16#0993# else
		x"852D" when address_in = 16#0994# else
		x"853E" when address_in = 16#0995# else
		x"2B23" when address_in = 16#0996# else
		x"F041" when address_in = 16#0997# else
		x"858F" when address_in = 16#0998# else
		x"8998" when address_in = 16#0999# else
		x"9595" when address_in = 16#099A# else
		x"9587" when address_in = 16#099B# else
		x"878F" when address_in = 16#099C# else
		x"8B98" when address_in = 16#099D# else
		x"9455" when address_in = 16#099E# else
		x"9447" when address_in = 16#099F# else
		x"88AD" when address_in = 16#09A0# else
		x"88BE" when address_in = 16#09A1# else
		x"14A6" when address_in = 16#09A2# else
		x"04B7" when address_in = 16#09A3# else
		x"F00C" when address_in = 16#09A4# else
		x"C0BA" when address_in = 16#09A5# else
		x"2CFD" when address_in = 16#09A6# else
		x"2CEC" when address_in = 16#09A7# else
		x"0CEE" when address_in = 16#09A8# else
		x"1CFF" when address_in = 16#09A9# else
		x"89EB" when address_in = 16#09AA# else
		x"89FC" when address_in = 16#09AB# else
		x"0EEE" when address_in = 16#09AC# else
		x"1EFF" when address_in = 16#09AD# else
		x"8529" when address_in = 16#09AE# else
		x"853A" when address_in = 16#09AF# else
		x"0F22" when address_in = 16#09B0# else
		x"1F33" when address_in = 16#09B1# else
		x"8B29" when address_in = 16#09B2# else
		x"8B3A" when address_in = 16#09B3# else
		x"8029" when address_in = 16#09B4# else
		x"803A" when address_in = 16#09B5# else
		x"0C2E" when address_in = 16#09B6# else
		x"1C3F" when address_in = 16#09B7# else
		x"2DF3" when address_in = 16#09B8# else
		x"2DE2" when address_in = 16#09B9# else
		x"8120" when address_in = 16#09BA# else
		x"8131" when address_in = 16#09BB# else
		x"858F" when address_in = 16#09BC# else
		x"8998" when address_in = 16#09BD# else
		x"2F73" when address_in = 16#09BE# else
		x"2F62" when address_in = 16#09BF# else
		x"940E" when address_in = 16#09C0# else
		x"0B02" when address_in = 16#09C1# else
		x"0F99" when address_in = 16#09C2# else
		x"0B88" when address_in = 16#09C3# else
		x"0F99" when address_in = 16#09C4# else
		x"2F98" when address_in = 16#09C5# else
		x"1F88" when address_in = 16#09C6# else
		x"2F08" when address_in = 16#09C7# else
		x"2F19" when address_in = 16#09C8# else
		x"9515" when address_in = 16#09C9# else
		x"9507" when address_in = 16#09CA# else
		x"7081" when address_in = 16#09CB# else
		x"7090" when address_in = 16#09CC# else
		x"0F08" when address_in = 16#09CD# else
		x"1F19" when address_in = 16#09CE# else
		x"808B" when address_in = 16#09CF# else
		x"809C" when address_in = 16#09D0# else
		x"0C8E" when address_in = 16#09D1# else
		x"1C9F" when address_in = 16#09D2# else
		x"2DF9" when address_in = 16#09D3# else
		x"2DE8" when address_in = 16#09D4# else
		x"8120" when address_in = 16#09D5# else
		x"8131" when address_in = 16#09D6# else
		x"2D95" when address_in = 16#09D7# else
		x"2D84" when address_in = 16#09D8# else
		x"2F73" when address_in = 16#09D9# else
		x"2F62" when address_in = 16#09DA# else
		x"940E" when address_in = 16#09DB# else
		x"0B02" when address_in = 16#09DC# else
		x"0F99" when address_in = 16#09DD# else
		x"0B88" when address_in = 16#09DE# else
		x"0F99" when address_in = 16#09DF# else
		x"2F98" when address_in = 16#09E0# else
		x"1F88" when address_in = 16#09E1# else
		x"2F28" when address_in = 16#09E2# else
		x"2F39" when address_in = 16#09E3# else
		x"9535" when address_in = 16#09E4# else
		x"9527" when address_in = 16#09E5# else
		x"7081" when address_in = 16#09E6# else
		x"7090" when address_in = 16#09E7# else
		x"0F28" when address_in = 16#09E8# else
		x"1F39" when address_in = 16#09E9# else
		x"1B02" when address_in = 16#09EA# else
		x"0B13" when address_in = 16#09EB# else
		x"8120" when address_in = 16#09EC# else
		x"8131" when address_in = 16#09ED# else
		x"858F" when address_in = 16#09EE# else
		x"8998" when address_in = 16#09EF# else
		x"2F73" when address_in = 16#09F0# else
		x"2F62" when address_in = 16#09F1# else
		x"940E" when address_in = 16#09F2# else
		x"0B02" when address_in = 16#09F3# else
		x"0F99" when address_in = 16#09F4# else
		x"0B88" when address_in = 16#09F5# else
		x"0F99" when address_in = 16#09F6# else
		x"2F98" when address_in = 16#09F7# else
		x"1F88" when address_in = 16#09F8# else
		x"2FB9" when address_in = 16#09F9# else
		x"2FA8" when address_in = 16#09FA# else
		x"95B5" when address_in = 16#09FB# else
		x"95A7" when address_in = 16#09FC# else
		x"7081" when address_in = 16#09FD# else
		x"7090" when address_in = 16#09FE# else
		x"0FA8" when address_in = 16#09FF# else
		x"1FB9" when address_in = 16#0A00# else
		x"2DF3" when address_in = 16#0A01# else
		x"2DE2" when address_in = 16#0A02# else
		x"8120" when address_in = 16#0A03# else
		x"8131" when address_in = 16#0A04# else
		x"2D95" when address_in = 16#0A05# else
		x"2D84" when address_in = 16#0A06# else
		x"2F73" when address_in = 16#0A07# else
		x"2F62" when address_in = 16#0A08# else
		x"940E" when address_in = 16#0A09# else
		x"0B02" when address_in = 16#0A0A# else
		x"0F99" when address_in = 16#0A0B# else
		x"0B88" when address_in = 16#0A0C# else
		x"0F99" when address_in = 16#0A0D# else
		x"2F98" when address_in = 16#0A0E# else
		x"1F88" when address_in = 16#0A0F# else
		x"2F28" when address_in = 16#0A10# else
		x"2F39" when address_in = 16#0A11# else
		x"9535" when address_in = 16#0A12# else
		x"9527" when address_in = 16#0A13# else
		x"7081" when address_in = 16#0A14# else
		x"7090" when address_in = 16#0A15# else
		x"0F28" when address_in = 16#0A16# else
		x"1F39" when address_in = 16#0A17# else
		x"0FA2" when address_in = 16#0A18# else
		x"1FB3" when address_in = 16#0A19# else
		x"2D9B" when address_in = 16#0A1A# else
		x"2D8A" when address_in = 16#0A1B# else
		x"0D8A" when address_in = 16#0A1C# else
		x"1D9B" when address_in = 16#0A1D# else
		x"8129" when address_in = 16#0A1E# else
		x"813A" when address_in = 16#0A1F# else
		x"0F28" when address_in = 16#0A20# else
		x"1F39" when address_in = 16#0A21# else
		x"8B2F" when address_in = 16#0A22# else
		x"8F38" when address_in = 16#0A23# else
		x"2FF3" when address_in = 16#0A24# else
		x"2FE2" when address_in = 16#0A25# else
		x"8120" when address_in = 16#0A26# else
		x"8131" when address_in = 16#0A27# else
		x"814B" when address_in = 16#0A28# else
		x"815C" when address_in = 16#0A29# else
		x"0F48" when address_in = 16#0A2A# else
		x"1F59" when address_in = 16#0A2B# else
		x"2FF5" when address_in = 16#0A2C# else
		x"2FE4" when address_in = 16#0A2D# else
		x"8160" when address_in = 16#0A2E# else
		x"8171" when address_in = 16#0A2F# else
		x"858D" when address_in = 16#0A30# else
		x"859E" when address_in = 16#0A31# else
		x"2B89" when address_in = 16#0A32# else
		x"F021" when address_in = 16#0A33# else
		x"9535" when address_in = 16#0A34# else
		x"9527" when address_in = 16#0A35# else
		x"9575" when address_in = 16#0A36# else
		x"9567" when address_in = 16#0A37# else
		x"2F93" when address_in = 16#0A38# else
		x"2F82" when address_in = 16#0A39# else
		x"1B80" when address_in = 16#0A3A# else
		x"0B91" when address_in = 16#0A3B# else
		x"2DF3" when address_in = 16#0A3C# else
		x"2DE2" when address_in = 16#0A3D# else
		x"8380" when address_in = 16#0A3E# else
		x"8391" when address_in = 16#0A3F# else
		x"2F97" when address_in = 16#0A40# else
		x"2F86" when address_in = 16#0A41# else
		x"1B8A" when address_in = 16#0A42# else
		x"0B9B" when address_in = 16#0A43# else
		x"2DF9" when address_in = 16#0A44# else
		x"2DE8" when address_in = 16#0A45# else
		x"8380" when address_in = 16#0A46# else
		x"8391" when address_in = 16#0A47# else
		x"0F20" when address_in = 16#0A48# else
		x"1F31" when address_in = 16#0A49# else
		x"89EF" when address_in = 16#0A4A# else
		x"8DF8" when address_in = 16#0A4B# else
		x"8320" when address_in = 16#0A4C# else
		x"8331" when address_in = 16#0A4D# else
		x"0F6A" when address_in = 16#0A4E# else
		x"1F7B" when address_in = 16#0A4F# else
		x"2FF5" when address_in = 16#0A50# else
		x"2FE4" when address_in = 16#0A51# else
		x"8360" when address_in = 16#0A52# else
		x"8371" when address_in = 16#0A53# else
		x"8529" when address_in = 16#0A54# else
		x"853A" when address_in = 16#0A55# else
		x"0EA2" when address_in = 16#0A56# else
		x"1EB3" when address_in = 16#0A57# else
		x"8989" when address_in = 16#0A58# else
		x"899A" when address_in = 16#0A59# else
		x"0EE8" when address_in = 16#0A5A# else
		x"1EF9" when address_in = 16#0A5B# else
		x"14A6" when address_in = 16#0A5C# else
		x"04B7" when address_in = 16#0A5D# else
		x"F40C" when address_in = 16#0A5E# else
		x"CF54" when address_in = 16#0A5F# else
		x"89ED" when address_in = 16#0A60# else
		x"89FE" when address_in = 16#0A61# else
		x"9631" when address_in = 16#0A62# else
		x"8BED" when address_in = 16#0A63# else
		x"8BFE" when address_in = 16#0A64# else
		x"892B" when address_in = 16#0A65# else
		x"893C" when address_in = 16#0A66# else
		x"5F2E" when address_in = 16#0A67# else
		x"4F3F" when address_in = 16#0A68# else
		x"8B2B" when address_in = 16#0A69# else
		x"8B3C" when address_in = 16#0A6A# else
		x"15EC" when address_in = 16#0A6B# else
		x"05FD" when address_in = 16#0A6C# else
		x"F40C" when address_in = 16#0A6D# else
		x"CEFB" when address_in = 16#0A6E# else
		x"818F" when address_in = 16#0A6F# else
		x"8598" when address_in = 16#0A70# else
		x"9701" when address_in = 16#0A71# else
		x"838F" when address_in = 16#0A72# else
		x"8798" when address_in = 16#0A73# else
		x"84C9" when address_in = 16#0A74# else
		x"84DA" when address_in = 16#0A75# else
		x"CE9B" when address_in = 16#0A76# else
		x"858B" when address_in = 16#0A77# else
		x"859C" when address_in = 16#0A78# else
		x"9668" when address_in = 16#0A79# else
		x"B60F" when address_in = 16#0A7A# else
		x"94F8" when address_in = 16#0A7B# else
		x"BFDE" when address_in = 16#0A7C# else
		x"BE0F" when address_in = 16#0A7D# else
		x"BFCD" when address_in = 16#0A7E# else
		x"91DF" when address_in = 16#0A7F# else
		x"91CF" when address_in = 16#0A80# else
		x"911F" when address_in = 16#0A81# else
		x"910F" when address_in = 16#0A82# else
		x"90FF" when address_in = 16#0A83# else
		x"90EF" when address_in = 16#0A84# else
		x"90DF" when address_in = 16#0A85# else
		x"90CF" when address_in = 16#0A86# else
		x"90BF" when address_in = 16#0A87# else
		x"90AF" when address_in = 16#0A88# else
		x"909F" when address_in = 16#0A89# else
		x"908F" when address_in = 16#0A8A# else
		x"907F" when address_in = 16#0A8B# else
		x"906F" when address_in = 16#0A8C# else
		x"905F" when address_in = 16#0A8D# else
		x"904F" when address_in = 16#0A8E# else
		x"903F" when address_in = 16#0A8F# else
		x"902F" when address_in = 16#0A90# else
		x"9508" when address_in = 16#0A91# else
		x"928F" when address_in = 16#0A92# else
		x"929F" when address_in = 16#0A93# else
		x"92AF" when address_in = 16#0A94# else
		x"92BF" when address_in = 16#0A95# else
		x"92CF" when address_in = 16#0A96# else
		x"92DF" when address_in = 16#0A97# else
		x"92EF" when address_in = 16#0A98# else
		x"92FF" when address_in = 16#0A99# else
		x"930F" when address_in = 16#0A9A# else
		x"931F" when address_in = 16#0A9B# else
		x"93CF" when address_in = 16#0A9C# else
		x"93DF" when address_in = 16#0A9D# else
		x"2EA8" when address_in = 16#0A9E# else
		x"2EB9" when address_in = 16#0A9F# else
		x"2EE6" when address_in = 16#0AA0# else
		x"2EF7" when address_in = 16#0AA1# else
		x"2EC4" when address_in = 16#0AA2# else
		x"2ED5" when address_in = 16#0AA3# else
		x"9408" when address_in = 16#0AA4# else
		x"08E1" when address_in = 16#0AA5# else
		x"08F1" when address_in = 16#0AA6# else
		x"E0A1" when address_in = 16#0AA7# else
		x"2E8A" when address_in = 16#0AA8# else
		x"2C91" when address_in = 16#0AA9# else
		x"2D19" when address_in = 16#0AAA# else
		x"2D08" when address_in = 16#0AAB# else
		x"2C0E" when address_in = 16#0AAC# else
		x"C002" when address_in = 16#0AAD# else
		x"0F00" when address_in = 16#0AAE# else
		x"1F11" when address_in = 16#0AAF# else
		x"940A" when address_in = 16#0AB0# else
		x"F7E2" when address_in = 16#0AB1# else
		x"E060" when address_in = 16#0AB2# else
		x"E070" when address_in = 16#0AB3# else
		x"2FD1" when address_in = 16#0AB4# else
		x"2FC0" when address_in = 16#0AB5# else
		x"0FC0" when address_in = 16#0AB6# else
		x"1FD1" when address_in = 16#0AB7# else
		x"0FC8" when address_in = 16#0AB8# else
		x"1FD9" when address_in = 16#0AB9# else
		x"1541" when address_in = 16#0ABA# else
		x"0551" when address_in = 16#0ABB# else
		x"F061" when address_in = 16#0ABC# else
		x"2F24" when address_in = 16#0ABD# else
		x"2F35" when address_in = 16#0ABE# else
		x"2D5F" when address_in = 16#0ABF# else
		x"2D4E" when address_in = 16#0AC0# else
		x"2F68" when address_in = 16#0AC1# else
		x"2F79" when address_in = 16#0AC2# else
		x"2F8C" when address_in = 16#0AC3# else
		x"2F9D" when address_in = 16#0AC4# else
		x"940E" when address_in = 16#0AC5# else
		x"0870" when address_in = 16#0AC6# else
		x"2F68" when address_in = 16#0AC7# else
		x"2F79" when address_in = 16#0AC8# else
		x"2D59" when address_in = 16#0AC9# else
		x"2D48" when address_in = 16#0ACA# else
		x"1680" when address_in = 16#0ACB# else
		x"0691" when address_in = 16#0ACC# else
		x"F4B4" when address_in = 16#0ACD# else
		x"2DBB" when address_in = 16#0ACE# else
		x"2DAA" when address_in = 16#0ACF# else
		x"9612" when address_in = 16#0AD0# else
		x"2FFD" when address_in = 16#0AD1# else
		x"2FEC" when address_in = 16#0AD2# else
		x"8120" when address_in = 16#0AD3# else
		x"8131" when address_in = 16#0AD4# else
		x"918D" when address_in = 16#0AD5# else
		x"919C" when address_in = 16#0AD6# else
		x"9711" when address_in = 16#0AD7# else
		x"8380" when address_in = 16#0AD8# else
		x"8391" when address_in = 16#0AD9# else
		x"932D" when address_in = 16#0ADA# else
		x"933C" when address_in = 16#0ADB# else
		x"9711" when address_in = 16#0ADC# else
		x"5F4E" when address_in = 16#0ADD# else
		x"4F5F" when address_in = 16#0ADE# else
		x"9634" when address_in = 16#0ADF# else
		x"9614" when address_in = 16#0AE0# else
		x"1740" when address_in = 16#0AE1# else
		x"0751" when address_in = 16#0AE2# else
		x"F37C" when address_in = 16#0AE3# else
		x"14C1" when address_in = 16#0AE4# else
		x"04D1" when address_in = 16#0AE5# else
		x"F461" when address_in = 16#0AE6# else
		x"2D3D" when address_in = 16#0AE7# else
		x"2D2C" when address_in = 16#0AE8# else
		x"2D5F" when address_in = 16#0AE9# else
		x"2D4E" when address_in = 16#0AEA# else
		x"2D7B" when address_in = 16#0AEB# else
		x"2D6A" when address_in = 16#0AEC# else
		x"2F8C" when address_in = 16#0AED# else
		x"2F9D" when address_in = 16#0AEE# else
		x"940E" when address_in = 16#0AEF# else
		x"0870" when address_in = 16#0AF0# else
		x"2F68" when address_in = 16#0AF1# else
		x"2F79" when address_in = 16#0AF2# else
		x"2F97" when address_in = 16#0AF3# else
		x"2F86" when address_in = 16#0AF4# else
		x"91DF" when address_in = 16#0AF5# else
		x"91CF" when address_in = 16#0AF6# else
		x"911F" when address_in = 16#0AF7# else
		x"910F" when address_in = 16#0AF8# else
		x"90FF" when address_in = 16#0AF9# else
		x"90EF" when address_in = 16#0AFA# else
		x"90DF" when address_in = 16#0AFB# else
		x"90CF" when address_in = 16#0AFC# else
		x"90BF" when address_in = 16#0AFD# else
		x"90AF" when address_in = 16#0AFE# else
		x"909F" when address_in = 16#0AFF# else
		x"908F" when address_in = 16#0B00# else
		x"9508" when address_in = 16#0B01# else
		x"2755" when address_in = 16#0B02# else
		x"2400" when address_in = 16#0B03# else
		x"FF80" when address_in = 16#0B04# else
		x"C002" when address_in = 16#0B05# else
		x"0E06" when address_in = 16#0B06# else
		x"1F57" when address_in = 16#0B07# else
		x"0F66" when address_in = 16#0B08# else
		x"1F77" when address_in = 16#0B09# else
		x"1561" when address_in = 16#0B0A# else
		x"0571" when address_in = 16#0B0B# else
		x"F021" when address_in = 16#0B0C# else
		x"9596" when address_in = 16#0B0D# else
		x"9587" when address_in = 16#0B0E# else
		x"9700" when address_in = 16#0B0F# else
		x"F799" when address_in = 16#0B10# else
		x"2F95" when address_in = 16#0B11# else
		x"2D80" when address_in = 16#0B12# else
		x"9508" when address_in = 16#0B13# else
		x"940C" when address_in = 16#1000# else
		x"0465" when address_in = 16#1001# else
		x"940C" when address_in = 16#1080# else
		x"0A92" when address_in = 16#1081# else
		x"940C" when address_in = 16#1380# else
		x"0565" when address_in = 16#1381# else
		x"940C" when address_in = 16#1382# else
		x"060F" when address_in = 16#1383# else
		x"940C" when address_in = 16#1384# else
		x"0692" when address_in = 16#1385# else
		x"ffff";
end rtl;
