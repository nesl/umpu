-- Input HEX file name : port_avr.ihex
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity programToLoad is port (
address_in : in  std_logic_vector (15 downto 0);
data_out   : out std_logic_vector (15 downto 0));
end programToLoad;

architecture rtl of programToLoad is
begin
data_out <=
		x"940C" when address_in = 16#0000# else
		x"0030" when address_in = 16#0001# else
		x"940C" when address_in = 16#0002# else
		x"0050" when address_in = 16#0003# else
		x"940C" when address_in = 16#0004# else
		x"0050" when address_in = 16#0005# else
		x"940C" when address_in = 16#0006# else
		x"0050" when address_in = 16#0007# else
		x"940C" when address_in = 16#0008# else
		x"0050" when address_in = 16#0009# else
		x"940C" when address_in = 16#000A# else
		x"0050" when address_in = 16#000B# else
		x"940C" when address_in = 16#000C# else
		x"0050" when address_in = 16#000D# else
		x"940C" when address_in = 16#000E# else
		x"0050" when address_in = 16#000F# else
		x"940C" when address_in = 16#0010# else
		x"0050" when address_in = 16#0011# else
		x"940C" when address_in = 16#0012# else
		x"0050" when address_in = 16#0013# else
		x"940C" when address_in = 16#0014# else
		x"0050" when address_in = 16#0015# else
		x"940C" when address_in = 16#0016# else
		x"0050" when address_in = 16#0017# else
		x"940C" when address_in = 16#0018# else
		x"0050" when address_in = 16#0019# else
		x"940C" when address_in = 16#001A# else
		x"0050" when address_in = 16#001B# else
		x"940C" when address_in = 16#001C# else
		x"0050" when address_in = 16#001D# else
		x"940C" when address_in = 16#001E# else
		x"00E9" when address_in = 16#001F# else
		x"940C" when address_in = 16#0020# else
		x"0050" when address_in = 16#0021# else
		x"940C" when address_in = 16#0022# else
		x"0050" when address_in = 16#0023# else
		x"940C" when address_in = 16#0024# else
		x"0050" when address_in = 16#0025# else
		x"940C" when address_in = 16#0026# else
		x"0050" when address_in = 16#0027# else
		x"940C" when address_in = 16#0028# else
		x"0050" when address_in = 16#0029# else
		x"940C" when address_in = 16#002A# else
		x"0050" when address_in = 16#002B# else
		x"940C" when address_in = 16#002C# else
		x"0050" when address_in = 16#002D# else
		x"940C" when address_in = 16#002E# else
		x"0050" when address_in = 16#002F# else
		x"2411" when address_in = 16#0030# else
		x"BE1F" when address_in = 16#0031# else
		x"EFCF" when address_in = 16#0032# else
		x"E0DF" when address_in = 16#0033# else
		x"BFDE" when address_in = 16#0034# else
		x"BFCD" when address_in = 16#0035# else
		x"E010" when address_in = 16#0036# else
		x"E6A0" when address_in = 16#0037# else
		x"E0B0" when address_in = 16#0038# else
		x"E9EA" when address_in = 16#0039# else
		x"E0F4" when address_in = 16#003A# else
		x"EF0F" when address_in = 16#003B# else
		x"9503" when address_in = 16#003C# else
		x"BF0B" when address_in = 16#003D# else
		x"C004" when address_in = 16#003E# else
		x"95D8" when address_in = 16#003F# else
		x"920D" when address_in = 16#0040# else
		x"9631" when address_in = 16#0041# else
		x"F3C8" when address_in = 16#0042# else
		x"36A0" when address_in = 16#0043# else
		x"07B1" when address_in = 16#0044# else
		x"F7C9" when address_in = 16#0045# else
		x"E010" when address_in = 16#0046# else
		x"E6A0" when address_in = 16#0047# else
		x"E0B0" when address_in = 16#0048# else
		x"C001" when address_in = 16#0049# else
		x"921D" when address_in = 16#004A# else
		x"38AD" when address_in = 16#004B# else
		x"07B1" when address_in = 16#004C# else
		x"F7E1" when address_in = 16#004D# else
		x"940C" when address_in = 16#004E# else
		x"0056" when address_in = 16#004F# else
		x"940C" when address_in = 16#0050# else
		x"0000" when address_in = 16#0051# else
		x"B38B" when address_in = 16#0052# else
		x"9580" when address_in = 16#0053# else
		x"BB8B" when address_in = 16#0054# else
		x"9508" when address_in = 16#0055# else
		x"EFCF" when address_in = 16#0056# else
		x"E0DF" when address_in = 16#0057# else
		x"BFDE" when address_in = 16#0058# else
		x"BFCD" when address_in = 16#0059# else
		x"940E" when address_in = 16#005A# else
		x"01EF" when address_in = 16#005B# else
		x"940E" when address_in = 16#005C# else
		x"01CD" when address_in = 16#005D# else
		x"9478" when address_in = 16#005E# else
		x"E522" when address_in = 16#005F# else
		x"E030" when address_in = 16#0060# else
		x"E644" when address_in = 16#0061# else
		x"E050" when address_in = 16#0062# else
		x"E16E" when address_in = 16#0063# else
		x"E070" when address_in = 16#0064# else
		x"E680" when address_in = 16#0065# else
		x"E090" when address_in = 16#0066# else
		x"940E" when address_in = 16#0067# else
		x"0184" when address_in = 16#0068# else
		x"EF8F" when address_in = 16#0069# else
		x"BB8A" when address_in = 16#006A# else
		x"BB8B" when address_in = 16#006B# else
		x"940E" when address_in = 16#006C# else
		x"021B" when address_in = 16#006D# else
		x"CFFF" when address_in = 16#006E# else
		x"93CF" when address_in = 16#006F# else
		x"93DF" when address_in = 16#0070# else
		x"2FB9" when address_in = 16#0071# else
		x"2FA8" when address_in = 16#0072# else
		x"E0C0" when address_in = 16#0073# else
		x"E0D0" when address_in = 16#0074# else
		x"91E0" when address_in = 16#0075# else
		x"0068" when address_in = 16#0076# else
		x"91F0" when address_in = 16#0077# else
		x"0069" when address_in = 16#0078# else
		x"2F4E" when address_in = 16#0079# else
		x"2F5F" when address_in = 16#007A# else
		x"9730" when address_in = 16#007B# else
		x"F0B1" when address_in = 16#007C# else
		x"8120" when address_in = 16#007D# else
		x"8131" when address_in = 16#007E# else
		x"918D" when address_in = 16#007F# else
		x"919C" when address_in = 16#0080# else
		x"9711" when address_in = 16#0081# else
		x"1782" when address_in = 16#0082# else
		x"0793" when address_in = 16#0083# else
		x"F0B8" when address_in = 16#0084# else
		x"1B82" when address_in = 16#0085# else
		x"0B93" when address_in = 16#0086# else
		x"938D" when address_in = 16#0087# else
		x"939C" when address_in = 16#0088# else
		x"9711" when address_in = 16#0089# else
		x"2FCE" when address_in = 16#008A# else
		x"2FDF" when address_in = 16#008B# else
		x"8006" when address_in = 16#008C# else
		x"81F7" when address_in = 16#008D# else
		x"2DE0" when address_in = 16#008E# else
		x"9730" when address_in = 16#008F# else
		x"F761" when address_in = 16#0090# else
		x"9720" when address_in = 16#0091# else
		x"F471" when address_in = 16#0092# else
		x"2FDB" when address_in = 16#0093# else
		x"2FCA" when address_in = 16#0094# else
		x"834E" when address_in = 16#0095# else
		x"835F" when address_in = 16#0096# else
		x"93B0" when address_in = 16#0097# else
		x"0069" when address_in = 16#0098# else
		x"93A0" when address_in = 16#0099# else
		x"0068" when address_in = 16#009A# else
		x"C00B" when address_in = 16#009B# else
		x"1B28" when address_in = 16#009C# else
		x"0B39" when address_in = 16#009D# else
		x"8320" when address_in = 16#009E# else
		x"8331" when address_in = 16#009F# else
		x"CFF0" when address_in = 16#00A0# else
		x"83AE" when address_in = 16#00A1# else
		x"83BF" when address_in = 16#00A2# else
		x"2FDB" when address_in = 16#00A3# else
		x"2FCA" when address_in = 16#00A4# else
		x"83EE" when address_in = 16#00A5# else
		x"83FF" when address_in = 16#00A6# else
		x"91DF" when address_in = 16#00A7# else
		x"91CF" when address_in = 16#00A8# else
		x"9508" when address_in = 16#00A9# else
		x"91E0" when address_in = 16#00AA# else
		x"0068" when address_in = 16#00AB# else
		x"91F0" when address_in = 16#00AC# else
		x"0069" when address_in = 16#00AD# else
		x"9730" when address_in = 16#00AE# else
		x"F439" when address_in = 16#00AF# else
		x"B780" when address_in = 16#00B0# else
		x"2799" when address_in = 16#00B1# else
		x"7086" when address_in = 16#00B2# else
		x"7090" when address_in = 16#00B3# else
		x"2B89" when address_in = 16#00B4# else
		x"F7D1" when address_in = 16#00B5# else
		x"C022" when address_in = 16#00B6# else
		x"B606" when address_in = 16#00B7# else
		x"FC01" when address_in = 16#00B8# else
		x"C02D" when address_in = 16#00B9# else
		x"B782" when address_in = 16#00BA# else
		x"2799" when address_in = 16#00BB# else
		x"8120" when address_in = 16#00BC# else
		x"8131" when address_in = 16#00BD# else
		x"1728" when address_in = 16#00BE# else
		x"0739" when address_in = 16#00BF# else
		x"F018" when address_in = 16#00C0# else
		x"1521" when address_in = 16#00C1# else
		x"0531" when address_in = 16#00C2# else
		x"F429" when address_in = 16#00C3# else
		x"E081" when address_in = 16#00C4# else
		x"E090" when address_in = 16#00C5# else
		x"8380" when address_in = 16#00C6# else
		x"8391" when address_in = 16#00C7# else
		x"C004" when address_in = 16#00C8# else
		x"1B28" when address_in = 16#00C9# else
		x"0B39" when address_in = 16#00CA# else
		x"8320" when address_in = 16#00CB# else
		x"8331" when address_in = 16#00CC# else
		x"8180" when address_in = 16#00CD# else
		x"8191" when address_in = 16#00CE# else
		x"3F8F" when address_in = 16#00CF# else
		x"0591" when address_in = 16#00D0# else
		x"F059" when address_in = 16#00D1# else
		x"F050" when address_in = 16#00D2# else
		x"B780" when address_in = 16#00D3# else
		x"2799" when address_in = 16#00D4# else
		x"7086" when address_in = 16#00D5# else
		x"7090" when address_in = 16#00D6# else
		x"2B89" when address_in = 16#00D7# else
		x"F7D1" when address_in = 16#00D8# else
		x"BE12" when address_in = 16#00D9# else
		x"EF8E" when address_in = 16#00DA# else
		x"BF81" when address_in = 16#00DB# else
		x"9508" when address_in = 16#00DC# else
		x"B780" when address_in = 16#00DD# else
		x"2799" when address_in = 16#00DE# else
		x"7086" when address_in = 16#00DF# else
		x"7090" when address_in = 16#00E0# else
		x"2B89" when address_in = 16#00E1# else
		x"F7D1" when address_in = 16#00E2# else
		x"BE12" when address_in = 16#00E3# else
		x"8180" when address_in = 16#00E4# else
		x"5081" when address_in = 16#00E5# else
		x"BF81" when address_in = 16#00E6# else
		x"9508" when address_in = 16#00E7# else
		x"9508" when address_in = 16#00E8# else
		x"921F" when address_in = 16#00E9# else
		x"920F" when address_in = 16#00EA# else
		x"B60F" when address_in = 16#00EB# else
		x"920F" when address_in = 16#00EC# else
		x"2411" when address_in = 16#00ED# else
		x"932F" when address_in = 16#00EE# else
		x"933F" when address_in = 16#00EF# else
		x"934F" when address_in = 16#00F0# else
		x"935F" when address_in = 16#00F1# else
		x"936F" when address_in = 16#00F2# else
		x"937F" when address_in = 16#00F3# else
		x"938F" when address_in = 16#00F4# else
		x"939F" when address_in = 16#00F5# else
		x"93AF" when address_in = 16#00F6# else
		x"93BF" when address_in = 16#00F7# else
		x"93CF" when address_in = 16#00F8# else
		x"93DF" when address_in = 16#00F9# else
		x"93EF" when address_in = 16#00FA# else
		x"93FF" when address_in = 16#00FB# else
		x"9160" when address_in = 16#00FC# else
		x"0068" when address_in = 16#00FD# else
		x"9170" when address_in = 16#00FE# else
		x"0069" when address_in = 16#00FF# else
		x"1561" when address_in = 16#0100# else
		x"0571" when address_in = 16#0101# else
		x"F409" when address_in = 16#0102# else
		x"C03E" when address_in = 16#0103# else
		x"2FF7" when address_in = 16#0104# else
		x"2FE6" when address_in = 16#0105# else
		x"B781" when address_in = 16#0106# else
		x"2F48" when address_in = 16#0107# else
		x"2755" when address_in = 16#0108# else
		x"5F4F" when address_in = 16#0109# else
		x"4F5F" when address_in = 16#010A# else
		x"8120" when address_in = 16#010B# else
		x"8131" when address_in = 16#010C# else
		x"1724" when address_in = 16#010D# else
		x"0735" when address_in = 16#010E# else
		x"F028" when address_in = 16#010F# else
		x"1B24" when address_in = 16#0110# else
		x"0B35" when address_in = 16#0111# else
		x"8320" when address_in = 16#0112# else
		x"8331" when address_in = 16#0113# else
		x"C009" when address_in = 16#0114# else
		x"1B42" when address_in = 16#0115# else
		x"0B53" when address_in = 16#0116# else
		x"8210" when address_in = 16#0117# else
		x"8211" when address_in = 16#0118# else
		x"8006" when address_in = 16#0119# else
		x"81F7" when address_in = 16#011A# else
		x"2DE0" when address_in = 16#011B# else
		x"9730" when address_in = 16#011C# else
		x"F769" when address_in = 16#011D# else
		x"2FD7" when address_in = 16#011E# else
		x"2FC6" when address_in = 16#011F# else
		x"C01C" when address_in = 16#0120# else
		x"8188" when address_in = 16#0121# else
		x"8199" when address_in = 16#0122# else
		x"2B89" when address_in = 16#0123# else
		x"F4D1" when address_in = 16#0124# else
		x"818E" when address_in = 16#0125# else
		x"819F" when address_in = 16#0126# else
		x"9390" when address_in = 16#0127# else
		x"0069" when address_in = 16#0128# else
		x"9380" when address_in = 16#0129# else
		x"0068" when address_in = 16#012A# else
		x"818C" when address_in = 16#012B# else
		x"819D" when address_in = 16#012C# else
		x"940E" when address_in = 16#012D# else
		x"01FE" when address_in = 16#012E# else
		x"818A" when address_in = 16#012F# else
		x"819B" when address_in = 16#0130# else
		x"9700" when address_in = 16#0131# else
		x"F031" when address_in = 16#0132# else
		x"8388" when address_in = 16#0133# else
		x"8399" when address_in = 16#0134# else
		x"2F8C" when address_in = 16#0135# else
		x"2F9D" when address_in = 16#0136# else
		x"940E" when address_in = 16#0137# else
		x"006F" when address_in = 16#0138# else
		x"91C0" when address_in = 16#0139# else
		x"0068" when address_in = 16#013A# else
		x"91D0" when address_in = 16#013B# else
		x"0069" when address_in = 16#013C# else
		x"9720" when address_in = 16#013D# else
		x"F711" when address_in = 16#013E# else
		x"940E" when address_in = 16#013F# else
		x"00AA" when address_in = 16#0140# else
		x"0000" when address_in = 16#0141# else
		x"91FF" when address_in = 16#0142# else
		x"91EF" when address_in = 16#0143# else
		x"91DF" when address_in = 16#0144# else
		x"91CF" when address_in = 16#0145# else
		x"91BF" when address_in = 16#0146# else
		x"91AF" when address_in = 16#0147# else
		x"919F" when address_in = 16#0148# else
		x"918F" when address_in = 16#0149# else
		x"917F" when address_in = 16#014A# else
		x"916F" when address_in = 16#014B# else
		x"915F" when address_in = 16#014C# else
		x"914F" when address_in = 16#014D# else
		x"913F" when address_in = 16#014E# else
		x"912F" when address_in = 16#014F# else
		x"900F" when address_in = 16#0150# else
		x"BE0F" when address_in = 16#0151# else
		x"900F" when address_in = 16#0152# else
		x"901F" when address_in = 16#0153# else
		x"9518" when address_in = 16#0154# else
		x"93CF" when address_in = 16#0155# else
		x"93DF" when address_in = 16#0156# else
		x"E0C0" when address_in = 16#0157# else
		x"E0D0" when address_in = 16#0158# else
		x"91E0" when address_in = 16#0159# else
		x"0068" when address_in = 16#015A# else
		x"91F0" when address_in = 16#015B# else
		x"0069" when address_in = 16#015C# else
		x"9730" when address_in = 16#015D# else
		x"F101" when address_in = 16#015E# else
		x"81A6" when address_in = 16#015F# else
		x"81B7" when address_in = 16#0160# else
		x"17E8" when address_in = 16#0161# else
		x"07F9" when address_in = 16#0162# else
		x"F4B1" when address_in = 16#0163# else
		x"9710" when address_in = 16#0164# else
		x"F051" when address_in = 16#0165# else
		x"918D" when address_in = 16#0166# else
		x"919C" when address_in = 16#0167# else
		x"9711" when address_in = 16#0168# else
		x"8120" when address_in = 16#0169# else
		x"8131" when address_in = 16#016A# else
		x"0F82" when address_in = 16#016B# else
		x"1F93" when address_in = 16#016C# else
		x"938D" when address_in = 16#016D# else
		x"939C" when address_in = 16#016E# else
		x"9711" when address_in = 16#016F# else
		x"9720" when address_in = 16#0170# else
		x"F019" when address_in = 16#0171# else
		x"83AE" when address_in = 16#0172# else
		x"83BF" when address_in = 16#0173# else
		x"C00A" when address_in = 16#0174# else
		x"93B0" when address_in = 16#0175# else
		x"0069" when address_in = 16#0176# else
		x"93A0" when address_in = 16#0177# else
		x"0068" when address_in = 16#0178# else
		x"C005" when address_in = 16#0179# else
		x"2FCE" when address_in = 16#017A# else
		x"2FDF" when address_in = 16#017B# else
		x"2FFB" when address_in = 16#017C# else
		x"2FEA" when address_in = 16#017D# else
		x"CFDE" when address_in = 16#017E# else
		x"2F8E" when address_in = 16#017F# else
		x"2F9F" when address_in = 16#0180# else
		x"91DF" when address_in = 16#0181# else
		x"91CF" when address_in = 16#0182# else
		x"9508" when address_in = 16#0183# else
		x"92AF" when address_in = 16#0184# else
		x"92BF" when address_in = 16#0185# else
		x"92CF" when address_in = 16#0186# else
		x"92DF" when address_in = 16#0187# else
		x"92EF" when address_in = 16#0188# else
		x"92FF" when address_in = 16#0189# else
		x"930F" when address_in = 16#018A# else
		x"931F" when address_in = 16#018B# else
		x"93CF" when address_in = 16#018C# else
		x"2F08" when address_in = 16#018D# else
		x"2F19" when address_in = 16#018E# else
		x"2EE6" when address_in = 16#018F# else
		x"2EF7" when address_in = 16#0190# else
		x"2EC4" when address_in = 16#0191# else
		x"2ED5" when address_in = 16#0192# else
		x"2EA2" when address_in = 16#0193# else
		x"2EB3" when address_in = 16#0194# else
		x"B7CF" when address_in = 16#0195# else
		x"94F8" when address_in = 16#0196# else
		x"940E" when address_in = 16#0197# else
		x"0155" when address_in = 16#0198# else
		x"2FF1" when address_in = 16#0199# else
		x"2FE0" when address_in = 16#019A# else
		x"82E0" when address_in = 16#019B# else
		x"82F1" when address_in = 16#019C# else
		x"82C2" when address_in = 16#019D# else
		x"82D3" when address_in = 16#019E# else
		x"82A4" when address_in = 16#019F# else
		x"82B5" when address_in = 16#01A0# else
		x"8216" when address_in = 16#01A1# else
		x"8217" when address_in = 16#01A2# else
		x"B782" when address_in = 16#01A3# else
		x"0EE8" when address_in = 16#01A4# else
		x"1CF1" when address_in = 16#01A5# else
		x"82E0" when address_in = 16#01A6# else
		x"82F1" when address_in = 16#01A7# else
		x"2F91" when address_in = 16#01A8# else
		x"2F80" when address_in = 16#01A9# else
		x"940E" when address_in = 16#01AA# else
		x"006F" when address_in = 16#01AB# else
		x"BFCF" when address_in = 16#01AC# else
		x"B7CF" when address_in = 16#01AD# else
		x"94F8" when address_in = 16#01AE# else
		x"940E" when address_in = 16#01AF# else
		x"00AA" when address_in = 16#01B0# else
		x"BFCF" when address_in = 16#01B1# else
		x"91CF" when address_in = 16#01B2# else
		x"911F" when address_in = 16#01B3# else
		x"910F" when address_in = 16#01B4# else
		x"90FF" when address_in = 16#01B5# else
		x"90EF" when address_in = 16#01B6# else
		x"90DF" when address_in = 16#01B7# else
		x"90CF" when address_in = 16#01B8# else
		x"90BF" when address_in = 16#01B9# else
		x"90AF" when address_in = 16#01BA# else
		x"9508" when address_in = 16#01BB# else
		x"93CF" when address_in = 16#01BC# else
		x"B7CF" when address_in = 16#01BD# else
		x"94F8" when address_in = 16#01BE# else
		x"940E" when address_in = 16#01BF# else
		x"0155" when address_in = 16#01C0# else
		x"2B89" when address_in = 16#01C1# else
		x"F039" when address_in = 16#01C2# else
		x"BFCF" when address_in = 16#01C3# else
		x"B7CF" when address_in = 16#01C4# else
		x"94F8" when address_in = 16#01C5# else
		x"940E" when address_in = 16#01C6# else
		x"00AA" when address_in = 16#01C7# else
		x"BFCF" when address_in = 16#01C8# else
		x"C001" when address_in = 16#01C9# else
		x"BFCF" when address_in = 16#01CA# else
		x"91CF" when address_in = 16#01CB# else
		x"9508" when address_in = 16#01CC# else
		x"9210" when address_in = 16#01CD# else
		x"0069" when address_in = 16#01CE# else
		x"9210" when address_in = 16#01CF# else
		x"0068" when address_in = 16#01D0# else
		x"940E" when address_in = 16#01D1# else
		x"01DD" when address_in = 16#01D2# else
		x"B780" when address_in = 16#01D3# else
		x"2799" when address_in = 16#01D4# else
		x"7086" when address_in = 16#01D5# else
		x"7090" when address_in = 16#01D6# else
		x"2B89" when address_in = 16#01D7# else
		x"F7D1" when address_in = 16#01D8# else
		x"BE12" when address_in = 16#01D9# else
		x"EF8E" when address_in = 16#01DA# else
		x"BF81" when address_in = 16#01DB# else
		x"9508" when address_in = 16#01DC# else
		x"B787" when address_in = 16#01DD# else
		x"7F8E" when address_in = 16#01DE# else
		x"BF87" when address_in = 16#01DF# else
		x"B787" when address_in = 16#01E0# else
		x"7F8D" when address_in = 16#01E1# else
		x"BF87" when address_in = 16#01E2# else
		x"B780" when address_in = 16#01E3# else
		x"6088" when address_in = 16#01E4# else
		x"BF80" when address_in = 16#01E5# else
		x"E089" when address_in = 16#01E6# else
		x"BF83" when address_in = 16#01E7# else
		x"BE12" when address_in = 16#01E8# else
		x"EF8F" when address_in = 16#01E9# else
		x"BF81" when address_in = 16#01EA# else
		x"B787" when address_in = 16#01EB# else
		x"6082" when address_in = 16#01EC# else
		x"BF87" when address_in = 16#01ED# else
		x"9508" when address_in = 16#01EE# else
		x"9210" when address_in = 16#01EF# else
		x"008A" when address_in = 16#01F0# else
		x"9210" when address_in = 16#01F1# else
		x"008B" when address_in = 16#01F2# else
		x"9210" when address_in = 16#01F3# else
		x"008C" when address_in = 16#01F4# else
		x"E08F" when address_in = 16#01F5# else
		x"E6EA" when address_in = 16#01F6# else
		x"E0F0" when address_in = 16#01F7# else
		x"9211" when address_in = 16#01F8# else
		x"9211" when address_in = 16#01F9# else
		x"5081" when address_in = 16#01FA# else
		x"FF87" when address_in = 16#01FB# else
		x"CFFB" when address_in = 16#01FC# else
		x"9508" when address_in = 16#01FD# else
		x"2F48" when address_in = 16#01FE# else
		x"2F59" when address_in = 16#01FF# else
		x"B73F" when address_in = 16#0200# else
		x"94F8" when address_in = 16#0201# else
		x"9120" when address_in = 16#0202# else
		x"008B" when address_in = 16#0203# else
		x"2FE2" when address_in = 16#0204# else
		x"27FF" when address_in = 16#0205# else
		x"0FEE" when address_in = 16#0206# else
		x"1FFF" when address_in = 16#0207# else
		x"59E6" when address_in = 16#0208# else
		x"4FFF" when address_in = 16#0209# else
		x"8180" when address_in = 16#020A# else
		x"8191" when address_in = 16#020B# else
		x"2B89" when address_in = 16#020C# else
		x"F459" when address_in = 16#020D# else
		x"5F2F" when address_in = 16#020E# else
		x"702F" when address_in = 16#020F# else
		x"9320" when address_in = 16#0210# else
		x"008B" when address_in = 16#0211# else
		x"8340" when address_in = 16#0212# else
		x"8351" when address_in = 16#0213# else
		x"9180" when address_in = 16#0214# else
		x"008C" when address_in = 16#0215# else
		x"5F8F" when address_in = 16#0216# else
		x"9380" when address_in = 16#0217# else
		x"008C" when address_in = 16#0218# else
		x"BF3F" when address_in = 16#0219# else
		x"9508" when address_in = 16#021A# else
		x"94F8" when address_in = 16#021B# else
		x"9180" when address_in = 16#021C# else
		x"008C" when address_in = 16#021D# else
		x"2388" when address_in = 16#021E# else
		x"F129" when address_in = 16#021F# else
		x"9478" when address_in = 16#0220# else
		x"9180" when address_in = 16#0221# else
		x"008A" when address_in = 16#0222# else
		x"2FE8" when address_in = 16#0223# else
		x"27FF" when address_in = 16#0224# else
		x"0FEE" when address_in = 16#0225# else
		x"1FFF" when address_in = 16#0226# else
		x"59E6" when address_in = 16#0227# else
		x"4FFF" when address_in = 16#0228# else
		x"8120" when address_in = 16#0229# else
		x"8131" when address_in = 16#022A# else
		x"9180" when address_in = 16#022B# else
		x"008A" when address_in = 16#022C# else
		x"2FE8" when address_in = 16#022D# else
		x"27FF" when address_in = 16#022E# else
		x"0FEE" when address_in = 16#022F# else
		x"1FFF" when address_in = 16#0230# else
		x"59E6" when address_in = 16#0231# else
		x"4FFF" when address_in = 16#0232# else
		x"8210" when address_in = 16#0233# else
		x"8211" when address_in = 16#0234# else
		x"9180" when address_in = 16#0235# else
		x"008A" when address_in = 16#0236# else
		x"5F8F" when address_in = 16#0237# else
		x"708F" when address_in = 16#0238# else
		x"9380" when address_in = 16#0239# else
		x"008A" when address_in = 16#023A# else
		x"9180" when address_in = 16#023B# else
		x"008C" when address_in = 16#023C# else
		x"5081" when address_in = 16#023D# else
		x"9380" when address_in = 16#023E# else
		x"008C" when address_in = 16#023F# else
		x"9478" when address_in = 16#0240# else
		x"2FE2" when address_in = 16#0241# else
		x"2FF3" when address_in = 16#0242# else
		x"9509" when address_in = 16#0243# else
		x"CFD6" when address_in = 16#0244# else
		x"B785" when address_in = 16#0245# else
		x"6280" when address_in = 16#0246# else
		x"BF85" when address_in = 16#0247# else
		x"9478" when address_in = 16#0248# else
		x"9588" when address_in = 16#0249# else
		x"0000" when address_in = 16#024A# else
		x"0000" when address_in = 16#024B# else
		x"CFCE" when address_in = 16#024C# else
		x"ffff";
end rtl;
