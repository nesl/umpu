-- Input HEX file name : test_mul_dom.ihex
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity programToLoad is port (
address_in : in  std_logic_vector (15 downto 0);
data_out   : out std_logic_vector (15 downto 0));
end programToLoad;

architecture rtl of programToLoad is
begin
data_out <=
		x"940C" when address_in = 16#0000# else
		x"0030" when address_in = 16#0001# else
		x"940C" when address_in = 16#0002# else
		x"0050" when address_in = 16#0003# else
		x"940C" when address_in = 16#0004# else
		x"0050" when address_in = 16#0005# else
		x"940C" when address_in = 16#0006# else
		x"0050" when address_in = 16#0007# else
		x"940C" when address_in = 16#0008# else
		x"0050" when address_in = 16#0009# else
		x"940C" when address_in = 16#000A# else
		x"0050" when address_in = 16#000B# else
		x"940C" when address_in = 16#000C# else
		x"0050" when address_in = 16#000D# else
		x"940C" when address_in = 16#000E# else
		x"0050" when address_in = 16#000F# else
		x"940C" when address_in = 16#0010# else
		x"0050" when address_in = 16#0011# else
		x"940C" when address_in = 16#0012# else
		x"0050" when address_in = 16#0013# else
		x"940C" when address_in = 16#0014# else
		x"0050" when address_in = 16#0015# else
		x"940C" when address_in = 16#0016# else
		x"0050" when address_in = 16#0017# else
		x"940C" when address_in = 16#0018# else
		x"0050" when address_in = 16#0019# else
		x"940C" when address_in = 16#001A# else
		x"0050" when address_in = 16#001B# else
		x"940C" when address_in = 16#001C# else
		x"0050" when address_in = 16#001D# else
		x"940C" when address_in = 16#001E# else
		x"0050" when address_in = 16#001F# else
		x"940C" when address_in = 16#0020# else
		x"0050" when address_in = 16#0021# else
		x"940C" when address_in = 16#0022# else
		x"0050" when address_in = 16#0023# else
		x"940C" when address_in = 16#0024# else
		x"0050" when address_in = 16#0025# else
		x"940C" when address_in = 16#0026# else
		x"0050" when address_in = 16#0027# else
		x"940C" when address_in = 16#0028# else
		x"0050" when address_in = 16#0029# else
		x"940C" when address_in = 16#002A# else
		x"00A1" when address_in = 16#002B# else
		x"940C" when address_in = 16#002C# else
		x"0050" when address_in = 16#002D# else
		x"940C" when address_in = 16#002E# else
		x"0050" when address_in = 16#002F# else
		x"2411" when address_in = 16#0030# else
		x"BE1F" when address_in = 16#0031# else
		x"EFCF" when address_in = 16#0032# else
		x"E0DF" when address_in = 16#0033# else
		x"BFDE" when address_in = 16#0034# else
		x"BFCD" when address_in = 16#0035# else
		x"E011" when address_in = 16#0036# else
		x"E6A0" when address_in = 16#0037# else
		x"E0B0" when address_in = 16#0038# else
		x"EBE6" when address_in = 16#0039# else
		x"E0F7" when address_in = 16#003A# else
		x"EF0F" when address_in = 16#003B# else
		x"9503" when address_in = 16#003C# else
		x"BF0B" when address_in = 16#003D# else
		x"C004" when address_in = 16#003E# else
		x"95D8" when address_in = 16#003F# else
		x"920D" when address_in = 16#0040# else
		x"9631" when address_in = 16#0041# else
		x"F3C8" when address_in = 16#0042# else
		x"36A0" when address_in = 16#0043# else
		x"07B1" when address_in = 16#0044# else
		x"F7C9" when address_in = 16#0045# else
		x"E011" when address_in = 16#0046# else
		x"E6A0" when address_in = 16#0047# else
		x"E0B1" when address_in = 16#0048# else
		x"C001" when address_in = 16#0049# else
		x"921D" when address_in = 16#004A# else
		x"36A6" when address_in = 16#004B# else
		x"07B1" when address_in = 16#004C# else
		x"F7E1" when address_in = 16#004D# else
		x"940C" when address_in = 16#004E# else
		x"0052" when address_in = 16#004F# else
		x"940C" when address_in = 16#0050# else
		x"0000" when address_in = 16#0051# else
		x"EFCF" when address_in = 16#0052# else
		x"E0DF" when address_in = 16#0053# else
		x"BFDE" when address_in = 16#0054# else
		x"BFCD" when address_in = 16#0055# else
		x"E688" when address_in = 16#0056# else
		x"B983" when address_in = 16#0057# else
		x"E089" when address_in = 16#0058# else
		x"B982" when address_in = 16#0059# else
		x"9478" when address_in = 16#005A# else
		x"940E" when address_in = 16#005B# else
		x"02A3" when address_in = 16#005C# else
		x"940E" when address_in = 16#005D# else
		x"1000" when address_in = 16#005E# else
		x"CFFF" when address_in = 16#005F# else
		x"2FF9" when address_in = 16#0060# else
		x"2FE8" when address_in = 16#0061# else
		x"E029" when address_in = 16#0062# else
		x"8180" when address_in = 16#0063# else
		x"2799" when address_in = 16#0064# else
		x"0F88" when address_in = 16#0065# else
		x"1F99" when address_in = 16#0066# else
		x"9381" when address_in = 16#0067# else
		x"BB8B" when address_in = 16#0068# else
		x"5021" when address_in = 16#0069# else
		x"FF27" when address_in = 16#006A# else
		x"CFF7" when address_in = 16#006B# else
		x"9508" when address_in = 16#006C# else
		x"93CF" when address_in = 16#006D# else
		x"93DF" when address_in = 16#006E# else
		x"EF8F" when address_in = 16#006F# else
		x"BB8A" when address_in = 16#0070# else
		x"B184" when address_in = 16#0071# else
		x"2799" when address_in = 16#0072# else
		x"718E" when address_in = 16#0073# else
		x"7090" when address_in = 16#0074# else
		x"9595" when address_in = 16#0075# else
		x"9587" when address_in = 16#0076# else
		x"9595" when address_in = 16#0077# else
		x"9587" when address_in = 16#0078# else
		x"2F68" when address_in = 16#0079# else
		x"E08A" when address_in = 16#007A# else
		x"E090" when address_in = 16#007B# else
		x"940E" when address_in = 16#007C# else
		x"1380" when address_in = 16#007D# else
		x"2FD9" when address_in = 16#007E# else
		x"2FC8" when address_in = 16#007F# else
		x"E080" when address_in = 16#0080# else
		x"2FFD" when address_in = 16#0081# else
		x"2FEC" when address_in = 16#0082# else
		x"9381" when address_in = 16#0083# else
		x"BB8B" when address_in = 16#0084# else
		x"5F8F" when address_in = 16#0085# else
		x"308A" when address_in = 16#0086# else
		x"F3D8" when address_in = 16#0087# else
		x"B184" when address_in = 16#0088# else
		x"2799" when address_in = 16#0089# else
		x"718E" when address_in = 16#008A# else
		x"7090" when address_in = 16#008B# else
		x"9595" when address_in = 16#008C# else
		x"9587" when address_in = 16#008D# else
		x"9595" when address_in = 16#008E# else
		x"9587" when address_in = 16#008F# else
		x"E041" when address_in = 16#0090# else
		x"2F68" when address_in = 16#0091# else
		x"2F8C" when address_in = 16#0092# else
		x"2F9D" when address_in = 16#0093# else
		x"940E" when address_in = 16#0094# else
		x"1384" when address_in = 16#0095# else
		x"2F8C" when address_in = 16#0096# else
		x"2F9D" when address_in = 16#0097# else
		x"940E" when address_in = 16#0098# else
		x"1080" when address_in = 16#0099# else
		x"E08A" when address_in = 16#009A# else
		x"8B8C" when address_in = 16#009B# else
		x"EF8F" when address_in = 16#009C# else
		x"BB8B" when address_in = 16#009D# else
		x"91DF" when address_in = 16#009E# else
		x"91CF" when address_in = 16#009F# else
		x"9508" when address_in = 16#00A0# else
		x"921F" when address_in = 16#00A1# else
		x"920F" when address_in = 16#00A2# else
		x"B60F" when address_in = 16#00A3# else
		x"920F" when address_in = 16#00A4# else
		x"2411" when address_in = 16#00A5# else
		x"938F" when address_in = 16#00A6# else
		x"E383" when address_in = 16#00A7# else
		x"BB8B" when address_in = 16#00A8# else
		x"EF80" when address_in = 16#00A9# else
		x"BB81" when address_in = 16#00AA# else
		x"E282" when address_in = 16#00AB# else
		x"BB8B" when address_in = 16#00AC# else
		x"CFFF" when address_in = 16#00AD# else
		x"93CF" when address_in = 16#00AE# else
		x"93DF" when address_in = 16#00AF# else
		x"2FF9" when address_in = 16#00B0# else
		x"2FE8" when address_in = 16#00B1# else
		x"81A2" when address_in = 16#00B2# else
		x"81B3" when address_in = 16#00B3# else
		x"8184" when address_in = 16#00B4# else
		x"8195" when address_in = 16#00B5# else
		x"2FDB" when address_in = 16#00B6# else
		x"2FCA" when address_in = 16#00B7# else
		x"838C" when address_in = 16#00B8# else
		x"839D" when address_in = 16#00B9# else
		x"8004" when address_in = 16#00BA# else
		x"81F5" when address_in = 16#00BB# else
		x"2DE0" when address_in = 16#00BC# else
		x"83A2" when address_in = 16#00BD# else
		x"83B3" when address_in = 16#00BE# else
		x"91DF" when address_in = 16#00BF# else
		x"91CF" when address_in = 16#00C0# else
		x"9508" when address_in = 16#00C1# else
		x"EF8F" when address_in = 16#00C2# else
		x"BB8B" when address_in = 16#00C3# else
		x"B38B" when address_in = 16#00C4# else
		x"9580" when address_in = 16#00C5# else
		x"CFFC" when address_in = 16#00C6# else
		x"93CF" when address_in = 16#00C7# else
		x"93DF" when address_in = 16#00C8# else
		x"2FF9" when address_in = 16#00C9# else
		x"2FE8" when address_in = 16#00CA# else
		x"91A0" when address_in = 16#00CB# else
		x"0162" when address_in = 16#00CC# else
		x"91B0" when address_in = 16#00CD# else
		x"0163" when address_in = 16#00CE# else
		x"2FDB" when address_in = 16#00CF# else
		x"2FCA" when address_in = 16#00D0# else
		x"818C" when address_in = 16#00D1# else
		x"819D" when address_in = 16#00D2# else
		x"83EC" when address_in = 16#00D3# else
		x"83FD" when address_in = 16#00D4# else
		x"83A2" when address_in = 16#00D5# else
		x"83B3" when address_in = 16#00D6# else
		x"8384" when address_in = 16#00D7# else
		x"8395" when address_in = 16#00D8# else
		x"2FD9" when address_in = 16#00D9# else
		x"2FC8" when address_in = 16#00DA# else
		x"83EA" when address_in = 16#00DB# else
		x"83FB" when address_in = 16#00DC# else
		x"91DF" when address_in = 16#00DD# else
		x"91CF" when address_in = 16#00DE# else
		x"9508" when address_in = 16#00DF# else
		x"92CF" when address_in = 16#00E0# else
		x"92DF" when address_in = 16#00E1# else
		x"92EF" when address_in = 16#00E2# else
		x"92FF" when address_in = 16#00E3# else
		x"930F" when address_in = 16#00E4# else
		x"931F" when address_in = 16#00E5# else
		x"93CF" when address_in = 16#00E6# else
		x"93DF" when address_in = 16#00E7# else
		x"2F16" when address_in = 16#00E8# else
		x"9700" when address_in = 16#00E9# else
		x"F409" when address_in = 16#00EA# else
		x"C095" when address_in = 16#00EB# else
		x"E059" when address_in = 16#00EC# else
		x"2EC5" when address_in = 16#00ED# else
		x"2CD1" when address_in = 16#00EE# else
		x"0EC8" when address_in = 16#00EF# else
		x"1ED9" when address_in = 16#00F0# else
		x"E043" when address_in = 16#00F1# else
		x"94D6" when address_in = 16#00F2# else
		x"94C7" when address_in = 16#00F3# else
		x"954A" when address_in = 16#00F4# else
		x"F7E1" when address_in = 16#00F5# else
		x"B70F" when address_in = 16#00F6# else
		x"94F8" when address_in = 16#00F7# else
		x"91E0" when address_in = 16#00F8# else
		x"0162" when address_in = 16#00F9# else
		x"91F0" when address_in = 16#00FA# else
		x"0163" when address_in = 16#00FB# else
		x"80E4" when address_in = 16#00FC# else
		x"80F5" when address_in = 16#00FD# else
		x"16EE" when address_in = 16#00FE# else
		x"06FF" when address_in = 16#00FF# else
		x"F181" when address_in = 16#0100# else
		x"2DBF" when address_in = 16#0101# else
		x"2DAE" when address_in = 16#0102# else
		x"91CD" when address_in = 16#0103# else
		x"91DC" when address_in = 16#0104# else
		x"E033" when address_in = 16#0105# else
		x"0FCC" when address_in = 16#0106# else
		x"1FDD" when address_in = 16#0107# else
		x"953A" when address_in = 16#0108# else
		x"F7E1" when address_in = 16#0109# else
		x"0DCE" when address_in = 16#010A# else
		x"1DDF" when address_in = 16#010B# else
		x"8188" when address_in = 16#010C# else
		x"8199" when address_in = 16#010D# else
		x"2399" when address_in = 16#010E# else
		x"F07C" when address_in = 16#010F# else
		x"2F8C" when address_in = 16#0110# else
		x"2F9D" when address_in = 16#0111# else
		x"940E" when address_in = 16#0112# else
		x"00AE" when address_in = 16#0113# else
		x"2DFF" when address_in = 16#0114# else
		x"2DEE" when address_in = 16#0115# else
		x"8180" when address_in = 16#0116# else
		x"8191" when address_in = 16#0117# else
		x"8128" when address_in = 16#0118# else
		x"8139" when address_in = 16#0119# else
		x"0F82" when address_in = 16#011A# else
		x"1F93" when address_in = 16#011B# else
		x"8380" when address_in = 16#011C# else
		x"8391" when address_in = 16#011D# else
		x"CFE2" when address_in = 16#011E# else
		x"2DBF" when address_in = 16#011F# else
		x"2DAE" when address_in = 16#0120# else
		x"918D" when address_in = 16#0121# else
		x"919C" when address_in = 16#0122# else
		x"158C" when address_in = 16#0123# else
		x"059D" when address_in = 16#0124# else
		x"F458" when address_in = 16#0125# else
		x"2DFF" when address_in = 16#0126# else
		x"2DEE" when address_in = 16#0127# else
		x"80E4" when address_in = 16#0128# else
		x"80F5" when address_in = 16#0129# else
		x"9180" when address_in = 16#012A# else
		x"0162" when address_in = 16#012B# else
		x"9190" when address_in = 16#012C# else
		x"0163" when address_in = 16#012D# else
		x"16E8" when address_in = 16#012E# else
		x"06F9" when address_in = 16#012F# else
		x"F681" when address_in = 16#0130# else
		x"9180" when address_in = 16#0131# else
		x"0162" when address_in = 16#0132# else
		x"9190" when address_in = 16#0133# else
		x"0163" when address_in = 16#0134# else
		x"16E8" when address_in = 16#0135# else
		x"06F9" when address_in = 16#0136# else
		x"F421" when address_in = 16#0137# else
		x"BF0F" when address_in = 16#0138# else
		x"E080" when address_in = 16#0139# else
		x"E090" when address_in = 16#013A# else
		x"C045" when address_in = 16#013B# else
		x"2DBF" when address_in = 16#013C# else
		x"2DAE" when address_in = 16#013D# else
		x"918D" when address_in = 16#013E# else
		x"919C" when address_in = 16#013F# else
		x"9711" when address_in = 16#0140# else
		x"16C8" when address_in = 16#0141# else
		x"06D9" when address_in = 16#0142# else
		x"F498" when address_in = 16#0143# else
		x"2DFD" when address_in = 16#0144# else
		x"2DEC" when address_in = 16#0145# else
		x"E023" when address_in = 16#0146# else
		x"0FEE" when address_in = 16#0147# else
		x"1FFF" when address_in = 16#0148# else
		x"952A" when address_in = 16#0149# else
		x"F7E1" when address_in = 16#014A# else
		x"0DEE" when address_in = 16#014B# else
		x"1DFF" when address_in = 16#014C# else
		x"198C" when address_in = 16#014D# else
		x"099D" when address_in = 16#014E# else
		x"8380" when address_in = 16#014F# else
		x"8391" when address_in = 16#0150# else
		x"92CD" when address_in = 16#0151# else
		x"92DC" when address_in = 16#0152# else
		x"2F8E" when address_in = 16#0153# else
		x"2F9F" when address_in = 16#0154# else
		x"940E" when address_in = 16#0155# else
		x"00C7" when address_in = 16#0156# else
		x"2D9F" when address_in = 16#0157# else
		x"2D8E" when address_in = 16#0158# else
		x"940E" when address_in = 16#0159# else
		x"00AE" when address_in = 16#015A# else
		x"2DFF" when address_in = 16#015B# else
		x"2DEE" when address_in = 16#015C# else
		x"8180" when address_in = 16#015D# else
		x"8191" when address_in = 16#015E# else
		x"6890" when address_in = 16#015F# else
		x"8380" when address_in = 16#0160# else
		x"8391" when address_in = 16#0161# else
		x"7017" when address_in = 16#0162# else
		x"2F81" when address_in = 16#0163# else
		x"6088" when address_in = 16#0164# else
		x"2F48" when address_in = 16#0165# else
		x"E068" when address_in = 16#0166# else
		x"E070" when address_in = 16#0167# else
		x"2D9F" when address_in = 16#0168# else
		x"2D8E" when address_in = 16#0169# else
		x"940E" when address_in = 16#016A# else
		x"0312" when address_in = 16#016B# else
		x"E083" when address_in = 16#016C# else
		x"0CCC" when address_in = 16#016D# else
		x"1CDD" when address_in = 16#016E# else
		x"958A" when address_in = 16#016F# else
		x"F7E1" when address_in = 16#0170# else
		x"EF88" when address_in = 16#0171# else
		x"EF9F" when address_in = 16#0172# else
		x"0EC8" when address_in = 16#0173# else
		x"1ED9" when address_in = 16#0174# else
		x"2F41" when address_in = 16#0175# else
		x"2D7D" when address_in = 16#0176# else
		x"2D6C" when address_in = 16#0177# else
		x"2D9F" when address_in = 16#0178# else
		x"2D8E" when address_in = 16#0179# else
		x"9608" when address_in = 16#017A# else
		x"940E" when address_in = 16#017B# else
		x"0312" when address_in = 16#017C# else
		x"BF0F" when address_in = 16#017D# else
		x"2D9F" when address_in = 16#017E# else
		x"2D8E" when address_in = 16#017F# else
		x"9602" when address_in = 16#0180# else
		x"91DF" when address_in = 16#0181# else
		x"91CF" when address_in = 16#0182# else
		x"911F" when address_in = 16#0183# else
		x"910F" when address_in = 16#0184# else
		x"90FF" when address_in = 16#0185# else
		x"90EF" when address_in = 16#0186# else
		x"90DF" when address_in = 16#0187# else
		x"90CF" when address_in = 16#0188# else
		x"9508" when address_in = 16#0189# else
		x"92EF" when address_in = 16#018A# else
		x"92FF" when address_in = 16#018B# else
		x"931F" when address_in = 16#018C# else
		x"93CF" when address_in = 16#018D# else
		x"93DF" when address_in = 16#018E# else
		x"2EE8" when address_in = 16#018F# else
		x"2EF9" when address_in = 16#0190# else
		x"9700" when address_in = 16#0191# else
		x"F409" when address_in = 16#0192# else
		x"C073" when address_in = 16#0193# else
		x"2FD9" when address_in = 16#0194# else
		x"2FC8" when address_in = 16#0195# else
		x"9722" when address_in = 16#0196# else
		x"E021" when address_in = 16#0197# else
		x"36C8" when address_in = 16#0198# else
		x"07D2" when address_in = 16#0199# else
		x"F408" when address_in = 16#019A# else
		x"C06B" when address_in = 16#019B# else
		x"9180" when address_in = 16#019C# else
		x"0164" when address_in = 16#019D# else
		x"9190" when address_in = 16#019E# else
		x"0165" when address_in = 16#019F# else
		x"E0A3" when address_in = 16#01A0# else
		x"0F88" when address_in = 16#01A1# else
		x"1F99" when address_in = 16#01A2# else
		x"95AA" when address_in = 16#01A3# else
		x"F7E1" when address_in = 16#01A4# else
		x"5988" when address_in = 16#01A5# else
		x"4F9E" when address_in = 16#01A6# else
		x"17C8" when address_in = 16#01A7# else
		x"07D9" when address_in = 16#01A8# else
		x"F008" when address_in = 16#01A9# else
		x"C05C" when address_in = 16#01AA# else
		x"B71F" when address_in = 16#01AB# else
		x"94F8" when address_in = 16#01AC# else
		x"B187" when address_in = 16#01AD# else
		x"2799" when address_in = 16#01AE# else
		x"2F98" when address_in = 16#01AF# else
		x"2788" when address_in = 16#01B0# else
		x"B128" when address_in = 16#01B1# else
		x"2733" when address_in = 16#01B2# else
		x"2B82" when address_in = 16#01B3# else
		x"2B93" when address_in = 16#01B4# else
		x"2F2C" when address_in = 16#01B5# else
		x"2F3D" when address_in = 16#01B6# else
		x"1B28" when address_in = 16#01B7# else
		x"0B39" when address_in = 16#01B8# else
		x"2FB3" when address_in = 16#01B9# else
		x"2FA2" when address_in = 16#01BA# else
		x"95B6" when address_in = 16#01BB# else
		x"95A7" when address_in = 16#01BC# else
		x"2FF3" when address_in = 16#01BD# else
		x"2FE2" when address_in = 16#01BE# else
		x"E074" when address_in = 16#01BF# else
		x"95F6" when address_in = 16#01C0# else
		x"95E7" when address_in = 16#01C1# else
		x"957A" when address_in = 16#01C2# else
		x"F7E1" when address_in = 16#01C3# else
		x"5AE0" when address_in = 16#01C4# else
		x"4FFF" when address_in = 16#01C5# else
		x"8140" when address_in = 16#01C6# else
		x"2F84" when address_in = 16#01C7# else
		x"2799" when address_in = 16#01C8# else
		x"70A4" when address_in = 16#01C9# else
		x"70B0" when address_in = 16#01CA# else
		x"2E0A" when address_in = 16#01CB# else
		x"C002" when address_in = 16#01CC# else
		x"9595" when address_in = 16#01CD# else
		x"9587" when address_in = 16#01CE# else
		x"940A" when address_in = 16#01CF# else
		x"F7E2" when address_in = 16#01D0# else
		x"2F48" when address_in = 16#01D1# else
		x"704F" when address_in = 16#01D2# else
		x"2F24" when address_in = 16#01D3# else
		x"2733" when address_in = 16#01D4# else
		x"2F93" when address_in = 16#01D5# else
		x"2F82" when address_in = 16#01D6# else
		x"7088" when address_in = 16#01D7# else
		x"7090" when address_in = 16#01D8# else
		x"5F87" when address_in = 16#01D9# else
		x"4F9F" when address_in = 16#01DA# else
		x"F411" when address_in = 16#01DB# else
		x"BF1F" when address_in = 16#01DC# else
		x"C008" when address_in = 16#01DD# else
		x"7027" when address_in = 16#01DE# else
		x"7030" when address_in = 16#01DF# else
		x"2F86" when address_in = 16#01E0# else
		x"2799" when address_in = 16#01E1# else
		x"1728" when address_in = 16#01E2# else
		x"0739" when address_in = 16#01E3# else
		x"F021" when address_in = 16#01E4# else
		x"BF1F" when address_in = 16#01E5# else
		x"940E" when address_in = 16#01E6# else
		x"00C2" when address_in = 16#01E7# else
		x"C01E" when address_in = 16#01E8# else
		x"B71F" when address_in = 16#01E9# else
		x"94F8" when address_in = 16#01EA# else
		x"8188" when address_in = 16#01EB# else
		x"8199" when address_in = 16#01EC# else
		x"779F" when address_in = 16#01ED# else
		x"8388" when address_in = 16#01EE# else
		x"8399" when address_in = 16#01EF# else
		x"8120" when address_in = 16#01F0# else
		x"E08F" when address_in = 16#01F1# else
		x"E090" when address_in = 16#01F2# else
		x"C002" when address_in = 16#01F3# else
		x"0F88" when address_in = 16#01F4# else
		x"1F99" when address_in = 16#01F5# else
		x"95AA" when address_in = 16#01F6# else
		x"F7E2" when address_in = 16#01F7# else
		x"2B28" when address_in = 16#01F8# else
		x"8320" when address_in = 16#01F9# else
		x"7047" when address_in = 16#01FA# else
		x"E02F" when address_in = 16#01FB# else
		x"2F62" when address_in = 16#01FC# else
		x"2D9F" when address_in = 16#01FD# else
		x"2D8E" when address_in = 16#01FE# else
		x"9606" when address_in = 16#01FF# else
		x"940E" when address_in = 16#0200# else
		x"036D" when address_in = 16#0201# else
		x"2F8C" when address_in = 16#0202# else
		x"2F9D" when address_in = 16#0203# else
		x"940E" when address_in = 16#0204# else
		x"00C7" when address_in = 16#0205# else
		x"BF1F" when address_in = 16#0206# else
		x"91DF" when address_in = 16#0207# else
		x"91CF" when address_in = 16#0208# else
		x"911F" when address_in = 16#0209# else
		x"90FF" when address_in = 16#020A# else
		x"90EF" when address_in = 16#020B# else
		x"9508" when address_in = 16#020C# else
		x"928F" when address_in = 16#020D# else
		x"929F" when address_in = 16#020E# else
		x"92AF" when address_in = 16#020F# else
		x"92BF" when address_in = 16#0210# else
		x"92CF" when address_in = 16#0211# else
		x"92DF" when address_in = 16#0212# else
		x"92EF" when address_in = 16#0213# else
		x"92FF" when address_in = 16#0214# else
		x"930F" when address_in = 16#0215# else
		x"931F" when address_in = 16#0216# else
		x"93CF" when address_in = 16#0217# else
		x"93DF" when address_in = 16#0218# else
		x"2EA8" when address_in = 16#0219# else
		x"2EB9" when address_in = 16#021A# else
		x"2E86" when address_in = 16#021B# else
		x"2E94" when address_in = 16#021C# else
		x"2F48" when address_in = 16#021D# else
		x"2F59" when address_in = 16#021E# else
		x"5042" when address_in = 16#021F# else
		x"4050" when address_in = 16#0220# else
		x"2B89" when address_in = 16#0221# else
		x"F409" when address_in = 16#0222# else
		x"C06C" when address_in = 16#0223# else
		x"B70F" when address_in = 16#0224# else
		x"94F8" when address_in = 16#0225# else
		x"B187" when address_in = 16#0226# else
		x"2799" when address_in = 16#0227# else
		x"2F98" when address_in = 16#0228# else
		x"2788" when address_in = 16#0229# else
		x"B128" when address_in = 16#022A# else
		x"2733" when address_in = 16#022B# else
		x"2B82" when address_in = 16#022C# else
		x"2B93" when address_in = 16#022D# else
		x"1B48" when address_in = 16#022E# else
		x"0B59" when address_in = 16#022F# else
		x"2EE4" when address_in = 16#0230# else
		x"2EF5" when address_in = 16#0231# else
		x"94F6" when address_in = 16#0232# else
		x"94E7" when address_in = 16#0233# else
		x"2EC4" when address_in = 16#0234# else
		x"2ED5" when address_in = 16#0235# else
		x"E0B4" when address_in = 16#0236# else
		x"94D6" when address_in = 16#0237# else
		x"94C7" when address_in = 16#0238# else
		x"95BA" when address_in = 16#0239# else
		x"F7E1" when address_in = 16#023A# else
		x"E680" when address_in = 16#023B# else
		x"E090" when address_in = 16#023C# else
		x"0EC8" when address_in = 16#023D# else
		x"1ED9" when address_in = 16#023E# else
		x"2DFD" when address_in = 16#023F# else
		x"2DEC" when address_in = 16#0240# else
		x"8110" when address_in = 16#0241# else
		x"2F81" when address_in = 16#0242# else
		x"2799" when address_in = 16#0243# else
		x"E0F4" when address_in = 16#0244# else
		x"22EF" when address_in = 16#0245# else
		x"24FF" when address_in = 16#0246# else
		x"2C0E" when address_in = 16#0247# else
		x"C002" when address_in = 16#0248# else
		x"9595" when address_in = 16#0249# else
		x"9587" when address_in = 16#024A# else
		x"940A" when address_in = 16#024B# else
		x"F7E2" when address_in = 16#024C# else
		x"2F18" when address_in = 16#024D# else
		x"701F" when address_in = 16#024E# else
		x"2FC1" when address_in = 16#024F# else
		x"27DD" when address_in = 16#0250# else
		x"2F8C" when address_in = 16#0251# else
		x"2F9D" when address_in = 16#0252# else
		x"7088" when address_in = 16#0253# else
		x"7090" when address_in = 16#0254# else
		x"5F87" when address_in = 16#0255# else
		x"4F9F" when address_in = 16#0256# else
		x"F419" when address_in = 16#0257# else
		x"BF0F" when address_in = 16#0258# else
		x"940E" when address_in = 16#0259# else
		x"00C2" when address_in = 16#025A# else
		x"2F2C" when address_in = 16#025B# else
		x"2F3D" when address_in = 16#025C# else
		x"7027" when address_in = 16#025D# else
		x"7030" when address_in = 16#025E# else
		x"2D88" when address_in = 16#025F# else
		x"2799" when address_in = 16#0260# else
		x"1728" when address_in = 16#0261# else
		x"0739" when address_in = 16#0262# else
		x"F549" when address_in = 16#0263# else
		x"2D49" when address_in = 16#0264# else
		x"2755" when address_in = 16#0265# else
		x"1742" when address_in = 16#0266# else
		x"0753" when address_in = 16#0267# else
		x"F151" when address_in = 16#0268# else
		x"2DFD" when address_in = 16#0269# else
		x"2DEC" when address_in = 16#026A# else
		x"8180" when address_in = 16#026B# else
		x"E02F" when address_in = 16#026C# else
		x"E030" when address_in = 16#026D# else
		x"2C0E" when address_in = 16#026E# else
		x"C002" when address_in = 16#026F# else
		x"0F22" when address_in = 16#0270# else
		x"1F33" when address_in = 16#0271# else
		x"940A" when address_in = 16#0272# else
		x"F7E2" when address_in = 16#0273# else
		x"2F92" when address_in = 16#0274# else
		x"9590" when address_in = 16#0275# else
		x"2389" when address_in = 16#0276# else
		x"7047" when address_in = 16#0277# else
		x"7050" when address_in = 16#0278# else
		x"6048" when address_in = 16#0279# else
		x"C002" when address_in = 16#027A# else
		x"0F44" when address_in = 16#027B# else
		x"1F55" when address_in = 16#027C# else
		x"94EA" when address_in = 16#027D# else
		x"F7E2" when address_in = 16#027E# else
		x"2B84" when address_in = 16#027F# else
		x"8380" when address_in = 16#0280# else
		x"E0F7" when address_in = 16#0281# else
		x"229F" when address_in = 16#0282# else
		x"231F" when address_in = 16#0283# else
		x"2D29" when address_in = 16#0284# else
		x"2F41" when address_in = 16#0285# else
		x"E06F" when address_in = 16#0286# else
		x"2D9B" when address_in = 16#0287# else
		x"2D8A" when address_in = 16#0288# else
		x"9606" when address_in = 16#0289# else
		x"940E" when address_in = 16#028A# else
		x"036D" when address_in = 16#028B# else
		x"C006" when address_in = 16#028C# else
		x"BF0F" when address_in = 16#028D# else
		x"940E" when address_in = 16#028E# else
		x"00C2" when address_in = 16#028F# else
		x"EF8F" when address_in = 16#0290# else
		x"EF9F" when address_in = 16#0291# else
		x"C003" when address_in = 16#0292# else
		x"BF0F" when address_in = 16#0293# else
		x"E080" when address_in = 16#0294# else
		x"E090" when address_in = 16#0295# else
		x"91DF" when address_in = 16#0296# else
		x"91CF" when address_in = 16#0297# else
		x"911F" when address_in = 16#0298# else
		x"910F" when address_in = 16#0299# else
		x"90FF" when address_in = 16#029A# else
		x"90EF" when address_in = 16#029B# else
		x"90DF" when address_in = 16#029C# else
		x"90CF" when address_in = 16#029D# else
		x"90BF" when address_in = 16#029E# else
		x"90AF" when address_in = 16#029F# else
		x"909F" when address_in = 16#02A0# else
		x"908F" when address_in = 16#02A1# else
		x"9508" when address_in = 16#02A2# else
		x"92EF" when address_in = 16#02A3# else
		x"92FF" when address_in = 16#02A4# else
		x"930F" when address_in = 16#02A5# else
		x"931F" when address_in = 16#02A6# else
		x"E608" when address_in = 16#02A7# else
		x"E011" when address_in = 16#02A8# else
		x"2CE1" when address_in = 16#02A9# else
		x"E038" when address_in = 16#02AA# else
		x"2EF3" when address_in = 16#02AB# else
		x"0EE0" when address_in = 16#02AC# else
		x"1EF1" when address_in = 16#02AD# else
		x"9310" when address_in = 16#02AE# else
		x"0161" when address_in = 16#02AF# else
		x"9300" when address_in = 16#02B0# else
		x"0160" when address_in = 16#02B1# else
		x"EF4F" when address_in = 16#02B2# else
		x"E050" when address_in = 16#02B3# else
		x"9350" when address_in = 16#02B4# else
		x"0165" when address_in = 16#02B5# else
		x"9340" when address_in = 16#02B6# else
		x"0164" when address_in = 16#02B7# else
		x"2F31" when address_in = 16#02B8# else
		x"2F20" when address_in = 16#02B9# else
		x"5028" when address_in = 16#02BA# else
		x"4F38" when address_in = 16#02BB# else
		x"9330" when address_in = 16#02BC# else
		x"0163" when address_in = 16#02BD# else
		x"9320" when address_in = 16#02BE# else
		x"0162" when address_in = 16#02BF# else
		x"E080" when address_in = 16#02C0# else
		x"E890" when address_in = 16#02C1# else
		x"9390" when address_in = 16#02C2# else
		x"0961" when address_in = 16#02C3# else
		x"9380" when address_in = 16#02C4# else
		x"0960" when address_in = 16#02C5# else
		x"9330" when address_in = 16#02C6# else
		x"0963" when address_in = 16#02C7# else
		x"9320" when address_in = 16#02C8# else
		x"0962" when address_in = 16#02C9# else
		x"9330" when address_in = 16#02CA# else
		x"0965" when address_in = 16#02CB# else
		x"9320" when address_in = 16#02CC# else
		x"0964" when address_in = 16#02CD# else
		x"9350" when address_in = 16#02CE# else
		x"0169" when address_in = 16#02CF# else
		x"9340" when address_in = 16#02D0# else
		x"0168" when address_in = 16#02D1# else
		x"2F91" when address_in = 16#02D2# else
		x"2F80" when address_in = 16#02D3# else
		x"940E" when address_in = 16#02D4# else
		x"00C7" when address_in = 16#02D5# else
		x"940E" when address_in = 16#02D6# else
		x"0308" when address_in = 16#02D7# else
		x"9180" when address_in = 16#02D8# else
		x"0164" when address_in = 16#02D9# else
		x"9190" when address_in = 16#02DA# else
		x"0165" when address_in = 16#02DB# else
		x"E023" when address_in = 16#02DC# else
		x"0F88" when address_in = 16#02DD# else
		x"1F99" when address_in = 16#02DE# else
		x"952A" when address_in = 16#02DF# else
		x"F7E1" when address_in = 16#02E0# else
		x"E04F" when address_in = 16#02E1# else
		x"2F68" when address_in = 16#02E2# else
		x"2F79" when address_in = 16#02E3# else
		x"9180" when address_in = 16#02E4# else
		x"0160" when address_in = 16#02E5# else
		x"9190" when address_in = 16#02E6# else
		x"0161" when address_in = 16#02E7# else
		x"940E" when address_in = 16#02E8# else
		x"0312" when address_in = 16#02E9# else
		x"B184" when address_in = 16#02EA# else
		x"718F" when address_in = 16#02EB# else
		x"B984" when address_in = 16#02EC# else
		x"B184" when address_in = 16#02ED# else
		x"6680" when address_in = 16#02EE# else
		x"B984" when address_in = 16#02EF# else
		x"9821" when address_in = 16#02F0# else
		x"B908" when address_in = 16#02F1# else
		x"2F81" when address_in = 16#02F2# else
		x"2799" when address_in = 16#02F3# else
		x"B987" when address_in = 16#02F4# else
		x"B8E6" when address_in = 16#02F5# else
		x"2D8F" when address_in = 16#02F6# else
		x"2799" when address_in = 16#02F7# else
		x"B985" when address_in = 16#02F8# else
		x"E680" when address_in = 16#02F9# else
		x"E090" when address_in = 16#02FA# else
		x"BB8D" when address_in = 16#02FB# else
		x"2F89" when address_in = 16#02FC# else
		x"2799" when address_in = 16#02FD# else
		x"BB8E" when address_in = 16#02FE# else
		x"BA1C" when address_in = 16#02FF# else
		x"E180" when address_in = 16#0300# else
		x"BB8F" when address_in = 16#0301# else
		x"9A20" when address_in = 16#0302# else
		x"911F" when address_in = 16#0303# else
		x"910F" when address_in = 16#0304# else
		x"90FF" when address_in = 16#0305# else
		x"90EF" when address_in = 16#0306# else
		x"9508" when address_in = 16#0307# else
		x"EF8F" when address_in = 16#0308# else
		x"E6E0" when address_in = 16#0309# else
		x"E0F0" when address_in = 16#030A# else
		x"9381" when address_in = 16#030B# else
		x"E091" when address_in = 16#030C# else
		x"35EF" when address_in = 16#030D# else
		x"07F9" when address_in = 16#030E# else
		x"F3D9" when address_in = 16#030F# else
		x"F3D0" when address_in = 16#0310# else
		x"9508" when address_in = 16#0311# else
		x"93CF" when address_in = 16#0312# else
		x"2FF9" when address_in = 16#0313# else
		x"2FE8" when address_in = 16#0314# else
		x"2FC4" when address_in = 16#0315# else
		x"1561" when address_in = 16#0316# else
		x"0571" when address_in = 16#0317# else
		x"F409" when address_in = 16#0318# else
		x"C051" when address_in = 16#0319# else
		x"2F97" when address_in = 16#031A# else
		x"2F86" when address_in = 16#031B# else
		x"7087" when address_in = 16#031C# else
		x"7F98" when address_in = 16#031D# else
		x"2B89" when address_in = 16#031E# else
		x"F009" when address_in = 16#031F# else
		x"C04A" when address_in = 16#0320# else
		x"E043" when address_in = 16#0321# else
		x"9576" when address_in = 16#0322# else
		x"9567" when address_in = 16#0323# else
		x"954A" when address_in = 16#0324# else
		x"F7E1" when address_in = 16#0325# else
		x"B187" when address_in = 16#0326# else
		x"2799" when address_in = 16#0327# else
		x"2F98" when address_in = 16#0328# else
		x"2788" when address_in = 16#0329# else
		x"B128" when address_in = 16#032A# else
		x"2733" when address_in = 16#032B# else
		x"2B82" when address_in = 16#032C# else
		x"2B93" when address_in = 16#032D# else
		x"1BE8" when address_in = 16#032E# else
		x"0BF9" when address_in = 16#032F# else
		x"2FAE" when address_in = 16#0330# else
		x"2FBF" when address_in = 16#0331# else
		x"E024" when address_in = 16#0332# else
		x"95B6" when address_in = 16#0333# else
		x"95A7" when address_in = 16#0334# else
		x"952A" when address_in = 16#0335# else
		x"F7E1" when address_in = 16#0336# else
		x"2F2E" when address_in = 16#0337# else
		x"2F3F" when address_in = 16#0338# else
		x"9536" when address_in = 16#0339# else
		x"9527" when address_in = 16#033A# else
		x"2FFB" when address_in = 16#033B# else
		x"2FEA" when address_in = 16#033C# else
		x"5AE0" when address_in = 16#033D# else
		x"4FFF" when address_in = 16#033E# else
		x"8150" when address_in = 16#033F# else
		x"7024" when address_in = 16#0340# else
		x"7030" when address_in = 16#0341# else
		x"E08F" when address_in = 16#0342# else
		x"E090" when address_in = 16#0343# else
		x"2E02" when address_in = 16#0344# else
		x"C002" when address_in = 16#0345# else
		x"0F88" when address_in = 16#0346# else
		x"1F99" when address_in = 16#0347# else
		x"940A" when address_in = 16#0348# else
		x"F7E2" when address_in = 16#0349# else
		x"2F48" when address_in = 16#034A# else
		x"2F8C" when address_in = 16#034B# else
		x"2799" when address_in = 16#034C# else
		x"C002" when address_in = 16#034D# else
		x"0F88" when address_in = 16#034E# else
		x"1F99" when address_in = 16#034F# else
		x"952A" when address_in = 16#0350# else
		x"F7E2" when address_in = 16#0351# else
		x"2F98" when address_in = 16#0352# else
		x"1561" when address_in = 16#0353# else
		x"0571" when address_in = 16#0354# else
		x"F091" when address_in = 16#0355# else
		x"2F84" when address_in = 16#0356# else
		x"9580" when address_in = 16#0357# else
		x"2358" when address_in = 16#0358# else
		x"2B59" when address_in = 16#0359# else
		x"5061" when address_in = 16#035A# else
		x"4070" when address_in = 16#035B# else
		x"9542" when address_in = 16#035C# else
		x"7F40" when address_in = 16#035D# else
		x"9592" when address_in = 16#035E# else
		x"7F90" when address_in = 16#035F# else
		x"2344" when address_in = 16#0360# else
		x"F789" when address_in = 16#0361# else
		x"9351" when address_in = 16#0362# else
		x"9611" when address_in = 16#0363# else
		x"8150" when address_in = 16#0364# else
		x"E04F" when address_in = 16#0365# else
		x"2F9C" when address_in = 16#0366# else
		x"CFEB" when address_in = 16#0367# else
		x"5AA0" when address_in = 16#0368# else
		x"4FBF" when address_in = 16#0369# else
		x"935C" when address_in = 16#036A# else
		x"91CF" when address_in = 16#036B# else
		x"9508" when address_in = 16#036C# else
		x"92FF" when address_in = 16#036D# else
		x"930F" when address_in = 16#036E# else
		x"931F" when address_in = 16#036F# else
		x"93CF" when address_in = 16#0370# else
		x"93DF" when address_in = 16#0371# else
		x"2EF6" when address_in = 16#0372# else
		x"2F04" when address_in = 16#0373# else
		x"2F12" when address_in = 16#0374# else
		x"E0C0" when address_in = 16#0375# else
		x"E0D0" when address_in = 16#0376# else
		x"B127" when address_in = 16#0377# else
		x"2733" when address_in = 16#0378# else
		x"2F32" when address_in = 16#0379# else
		x"2722" when address_in = 16#037A# else
		x"B148" when address_in = 16#037B# else
		x"2755" when address_in = 16#037C# else
		x"2B24" when address_in = 16#037D# else
		x"2B35" when address_in = 16#037E# else
		x"1B82" when address_in = 16#037F# else
		x"0B93" when address_in = 16#0380# else
		x"2FB9" when address_in = 16#0381# else
		x"2FA8" when address_in = 16#0382# else
		x"E064" when address_in = 16#0383# else
		x"95B6" when address_in = 16#0384# else
		x"95A7" when address_in = 16#0385# else
		x"956A" when address_in = 16#0386# else
		x"F7E1" when address_in = 16#0387# else
		x"2F28" when address_in = 16#0388# else
		x"2F39" when address_in = 16#0389# else
		x"9536" when address_in = 16#038A# else
		x"9527" when address_in = 16#038B# else
		x"2FFB" when address_in = 16#038C# else
		x"2FEA" when address_in = 16#038D# else
		x"5AE0" when address_in = 16#038E# else
		x"4FFF" when address_in = 16#038F# else
		x"8140" when address_in = 16#0390# else
		x"2D8F" when address_in = 16#0391# else
		x"2799" when address_in = 16#0392# else
		x"7024" when address_in = 16#0393# else
		x"7030" when address_in = 16#0394# else
		x"2E02" when address_in = 16#0395# else
		x"C002" when address_in = 16#0396# else
		x"0F88" when address_in = 16#0397# else
		x"1F99" when address_in = 16#0398# else
		x"940A" when address_in = 16#0399# else
		x"F7E2" when address_in = 16#039A# else
		x"2F68" when address_in = 16#039B# else
		x"2F80" when address_in = 16#039C# else
		x"2799" when address_in = 16#039D# else
		x"2E02" when address_in = 16#039E# else
		x"C002" when address_in = 16#039F# else
		x"0F88" when address_in = 16#03A0# else
		x"1F99" when address_in = 16#03A1# else
		x"940A" when address_in = 16#03A2# else
		x"F7E2" when address_in = 16#03A3# else
		x"2F58" when address_in = 16#03A4# else
		x"2F81" when address_in = 16#03A5# else
		x"2799" when address_in = 16#03A6# else
		x"2E02" when address_in = 16#03A7# else
		x"C002" when address_in = 16#03A8# else
		x"0F88" when address_in = 16#03A9# else
		x"1F99" when address_in = 16#03AA# else
		x"940A" when address_in = 16#03AB# else
		x"F7E2" when address_in = 16#03AC# else
		x"2F78" when address_in = 16#03AD# else
		x"E08F" when address_in = 16#03AE# else
		x"E090" when address_in = 16#03AF# else
		x"C002" when address_in = 16#03B0# else
		x"0F88" when address_in = 16#03B1# else
		x"1F99" when address_in = 16#03B2# else
		x"952A" when address_in = 16#03B3# else
		x"F7E2" when address_in = 16#03B4# else
		x"2F98" when address_in = 16#03B5# else
		x"2F84" when address_in = 16#03B6# else
		x"2386" when address_in = 16#03B7# else
		x"1785" when address_in = 16#03B8# else
		x"F4B1" when address_in = 16#03B9# else
		x"2F89" when address_in = 16#03BA# else
		x"9580" when address_in = 16#03BB# else
		x"2348" when address_in = 16#03BC# else
		x"2B47" when address_in = 16#03BD# else
		x"9621" when address_in = 16#03BE# else
		x"9562" when address_in = 16#03BF# else
		x"7F60" when address_in = 16#03C0# else
		x"9552" when address_in = 16#03C1# else
		x"7F50" when address_in = 16#03C2# else
		x"9572" when address_in = 16#03C3# else
		x"7F70" when address_in = 16#03C4# else
		x"9592" when address_in = 16#03C5# else
		x"7F90" when address_in = 16#03C6# else
		x"F771" when address_in = 16#03C7# else
		x"9341" when address_in = 16#03C8# else
		x"9611" when address_in = 16#03C9# else
		x"8140" when address_in = 16#03CA# else
		x"2D6F" when address_in = 16#03CB# else
		x"2F50" when address_in = 16#03CC# else
		x"2F71" when address_in = 16#03CD# else
		x"E09F" when address_in = 16#03CE# else
		x"CFE6" when address_in = 16#03CF# else
		x"5AA0" when address_in = 16#03D0# else
		x"4FBF" when address_in = 16#03D1# else
		x"934C" when address_in = 16#03D2# else
		x"2F8C" when address_in = 16#03D3# else
		x"2F9D" when address_in = 16#03D4# else
		x"91DF" when address_in = 16#03D5# else
		x"91CF" when address_in = 16#03D6# else
		x"911F" when address_in = 16#03D7# else
		x"910F" when address_in = 16#03D8# else
		x"90FF" when address_in = 16#03D9# else
		x"9508" when address_in = 16#03DA# else
		x"940C" when address_in = 16#1000# else
		x"006D" when address_in = 16#1001# else
		x"940C" when address_in = 16#1080# else
		x"0060" when address_in = 16#1081# else
		x"940C" when address_in = 16#1380# else
		x"00E0" when address_in = 16#1381# else
		x"940C" when address_in = 16#1382# else
		x"018A" when address_in = 16#1383# else
		x"940C" when address_in = 16#1384# else
		x"020D" when address_in = 16#1385# else
		x"ffff";
end rtl;
