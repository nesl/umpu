-- Input HEX file name : blink_app.ihex
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity programToLoad is port (
address_in : in  std_logic_vector (15 downto 0);
data_out   : out std_logic_vector (15 downto 0));
end programToLoad;

architecture rtl of programToLoad is
begin
data_out <=
		x"940C" when address_in = 16#0000# else
		x"0595" when address_in = 16#0001# else
		x"940C" when address_in = 16#0002# else
		x"05B5" when address_in = 16#0003# else
		x"940C" when address_in = 16#0004# else
		x"05B5" when address_in = 16#0005# else
		x"940C" when address_in = 16#0006# else
		x"05B5" when address_in = 16#0007# else
		x"940C" when address_in = 16#0008# else
		x"05B5" when address_in = 16#0009# else
		x"940C" when address_in = 16#000A# else
		x"05B5" when address_in = 16#000B# else
		x"940C" when address_in = 16#000C# else
		x"05B5" when address_in = 16#000D# else
		x"940C" when address_in = 16#000E# else
		x"05B5" when address_in = 16#000F# else
		x"940C" when address_in = 16#0010# else
		x"05B5" when address_in = 16#0011# else
		x"940C" when address_in = 16#0012# else
		x"05B5" when address_in = 16#0013# else
		x"940C" when address_in = 16#0014# else
		x"05B5" when address_in = 16#0015# else
		x"940C" when address_in = 16#0016# else
		x"05B5" when address_in = 16#0017# else
		x"940C" when address_in = 16#0018# else
		x"05B5" when address_in = 16#0019# else
		x"940C" when address_in = 16#001A# else
		x"05B5" when address_in = 16#001B# else
		x"940C" when address_in = 16#001C# else
		x"05B5" when address_in = 16#001D# else
		x"940C" when address_in = 16#001E# else
		x"2263" when address_in = 16#001F# else
		x"940C" when address_in = 16#0020# else
		x"05B5" when address_in = 16#0021# else
		x"940C" when address_in = 16#0022# else
		x"05B5" when address_in = 16#0023# else
		x"940C" when address_in = 16#0024# else
		x"29E4" when address_in = 16#0025# else
		x"940C" when address_in = 16#0026# else
		x"05B5" when address_in = 16#0027# else
		x"940C" when address_in = 16#0028# else
		x"27D2" when address_in = 16#0029# else
		x"940C" when address_in = 16#002A# else
		x"2E1F" when address_in = 16#002B# else
		x"940C" when address_in = 16#002C# else
		x"05B5" when address_in = 16#002D# else
		x"940C" when address_in = 16#002E# else
		x"05B5" when address_in = 16#002F# else
		x"0000" when address_in = 16#0030# else
		x"0000" when address_in = 16#0031# else
		x"0000" when address_in = 16#0032# else
		x"0000" when address_in = 16#0033# else
		x"0000" when address_in = 16#0034# else
		x"0000" when address_in = 16#0035# else
		x"0000" when address_in = 16#0036# else
		x"0000" when address_in = 16#0037# else
		x"0000" when address_in = 16#0038# else
		x"0000" when address_in = 16#0039# else
		x"0000" when address_in = 16#003A# else
		x"0000" when address_in = 16#003B# else
		x"0000" when address_in = 16#003C# else
		x"0000" when address_in = 16#003D# else
		x"0000" when address_in = 16#003E# else
		x"0000" when address_in = 16#003F# else
		x"0000" when address_in = 16#0040# else
		x"0000" when address_in = 16#0041# else
		x"0000" when address_in = 16#0042# else
		x"0000" when address_in = 16#0043# else
		x"0000" when address_in = 16#0044# else
		x"0000" when address_in = 16#0045# else
		x"0000" when address_in = 16#0046# else
		x"0000" when address_in = 16#0047# else
		x"0000" when address_in = 16#0048# else
		x"0000" when address_in = 16#0049# else
		x"0000" when address_in = 16#004A# else
		x"0000" when address_in = 16#004B# else
		x"0000" when address_in = 16#004C# else
		x"0000" when address_in = 16#004D# else
		x"0000" when address_in = 16#004E# else
		x"0000" when address_in = 16#004F# else
		x"0000" when address_in = 16#0050# else
		x"0000" when address_in = 16#0051# else
		x"0000" when address_in = 16#0052# else
		x"0000" when address_in = 16#0053# else
		x"0000" when address_in = 16#0054# else
		x"0000" when address_in = 16#0055# else
		x"0000" when address_in = 16#0056# else
		x"0000" when address_in = 16#0057# else
		x"0000" when address_in = 16#0058# else
		x"0000" when address_in = 16#0059# else
		x"0000" when address_in = 16#005A# else
		x"0000" when address_in = 16#005B# else
		x"0000" when address_in = 16#005C# else
		x"0000" when address_in = 16#005D# else
		x"0000" when address_in = 16#005E# else
		x"0000" when address_in = 16#005F# else
		x"0000" when address_in = 16#0060# else
		x"0000" when address_in = 16#0061# else
		x"0000" when address_in = 16#0062# else
		x"0000" when address_in = 16#0063# else
		x"0000" when address_in = 16#0064# else
		x"0000" when address_in = 16#0065# else
		x"0000" when address_in = 16#0066# else
		x"0000" when address_in = 16#0067# else
		x"0000" when address_in = 16#0068# else
		x"0000" when address_in = 16#0069# else
		x"0000" when address_in = 16#006A# else
		x"0000" when address_in = 16#006B# else
		x"0000" when address_in = 16#006C# else
		x"0000" when address_in = 16#006D# else
		x"0000" when address_in = 16#006E# else
		x"0000" when address_in = 16#006F# else
		x"0000" when address_in = 16#0070# else
		x"0000" when address_in = 16#0071# else
		x"0000" when address_in = 16#0072# else
		x"0000" when address_in = 16#0073# else
		x"0000" when address_in = 16#0074# else
		x"0000" when address_in = 16#0075# else
		x"0000" when address_in = 16#0076# else
		x"0000" when address_in = 16#0077# else
		x"0000" when address_in = 16#0078# else
		x"0000" when address_in = 16#0079# else
		x"0000" when address_in = 16#007A# else
		x"0000" when address_in = 16#007B# else
		x"0000" when address_in = 16#007C# else
		x"0000" when address_in = 16#007D# else
		x"0000" when address_in = 16#007E# else
		x"0000" when address_in = 16#007F# else
		x"940C" when address_in = 16#0080# else
		x"05F0" when address_in = 16#0081# else
		x"0000" when address_in = 16#0082# else
		x"0000" when address_in = 16#0083# else
		x"0000" when address_in = 16#0084# else
		x"0000" when address_in = 16#0085# else
		x"0000" when address_in = 16#0086# else
		x"0000" when address_in = 16#0087# else
		x"0000" when address_in = 16#0088# else
		x"0000" when address_in = 16#0089# else
		x"0000" when address_in = 16#008A# else
		x"0000" when address_in = 16#008B# else
		x"0000" when address_in = 16#008C# else
		x"0000" when address_in = 16#008D# else
		x"0000" when address_in = 16#008E# else
		x"0000" when address_in = 16#008F# else
		x"0000" when address_in = 16#0090# else
		x"0000" when address_in = 16#0091# else
		x"0000" when address_in = 16#0092# else
		x"0000" when address_in = 16#0093# else
		x"0000" when address_in = 16#0094# else
		x"0000" when address_in = 16#0095# else
		x"0000" when address_in = 16#0096# else
		x"0000" when address_in = 16#0097# else
		x"0000" when address_in = 16#0098# else
		x"0000" when address_in = 16#0099# else
		x"0000" when address_in = 16#009A# else
		x"0000" when address_in = 16#009B# else
		x"0000" when address_in = 16#009C# else
		x"0000" when address_in = 16#009D# else
		x"0000" when address_in = 16#009E# else
		x"0000" when address_in = 16#009F# else
		x"0000" when address_in = 16#00A0# else
		x"0000" when address_in = 16#00A1# else
		x"0000" when address_in = 16#00A2# else
		x"0000" when address_in = 16#00A3# else
		x"0000" when address_in = 16#00A4# else
		x"0000" when address_in = 16#00A5# else
		x"0000" when address_in = 16#00A6# else
		x"0000" when address_in = 16#00A7# else
		x"0000" when address_in = 16#00A8# else
		x"0000" when address_in = 16#00A9# else
		x"0000" when address_in = 16#00AA# else
		x"0000" when address_in = 16#00AB# else
		x"0000" when address_in = 16#00AC# else
		x"0000" when address_in = 16#00AD# else
		x"0000" when address_in = 16#00AE# else
		x"0000" when address_in = 16#00AF# else
		x"0000" when address_in = 16#00B0# else
		x"0000" when address_in = 16#00B1# else
		x"0000" when address_in = 16#00B2# else
		x"0000" when address_in = 16#00B3# else
		x"0000" when address_in = 16#00B4# else
		x"0000" when address_in = 16#00B5# else
		x"0000" when address_in = 16#00B6# else
		x"0000" when address_in = 16#00B7# else
		x"0000" when address_in = 16#00B8# else
		x"0000" when address_in = 16#00B9# else
		x"0000" when address_in = 16#00BA# else
		x"0000" when address_in = 16#00BB# else
		x"0000" when address_in = 16#00BC# else
		x"0000" when address_in = 16#00BD# else
		x"0000" when address_in = 16#00BE# else
		x"0000" when address_in = 16#00BF# else
		x"0000" when address_in = 16#00C0# else
		x"0000" when address_in = 16#00C1# else
		x"0000" when address_in = 16#00C2# else
		x"0000" when address_in = 16#00C3# else
		x"0000" when address_in = 16#00C4# else
		x"0000" when address_in = 16#00C5# else
		x"0000" when address_in = 16#00C6# else
		x"0000" when address_in = 16#00C7# else
		x"0000" when address_in = 16#00C8# else
		x"0000" when address_in = 16#00C9# else
		x"0000" when address_in = 16#00CA# else
		x"0000" when address_in = 16#00CB# else
		x"0000" when address_in = 16#00CC# else
		x"0000" when address_in = 16#00CD# else
		x"0000" when address_in = 16#00CE# else
		x"0000" when address_in = 16#00CF# else
		x"0000" when address_in = 16#00D0# else
		x"0000" when address_in = 16#00D1# else
		x"0000" when address_in = 16#00D2# else
		x"0000" when address_in = 16#00D3# else
		x"0000" when address_in = 16#00D4# else
		x"0000" when address_in = 16#00D5# else
		x"0000" when address_in = 16#00D6# else
		x"0000" when address_in = 16#00D7# else
		x"0000" when address_in = 16#00D8# else
		x"0000" when address_in = 16#00D9# else
		x"0000" when address_in = 16#00DA# else
		x"0000" when address_in = 16#00DB# else
		x"0000" when address_in = 16#00DC# else
		x"0000" when address_in = 16#00DD# else
		x"0000" when address_in = 16#00DE# else
		x"0000" when address_in = 16#00DF# else
		x"0000" when address_in = 16#00E0# else
		x"0000" when address_in = 16#00E1# else
		x"0000" when address_in = 16#00E2# else
		x"0000" when address_in = 16#00E3# else
		x"0000" when address_in = 16#00E4# else
		x"0000" when address_in = 16#00E5# else
		x"0000" when address_in = 16#00E6# else
		x"0000" when address_in = 16#00E7# else
		x"0000" when address_in = 16#00E8# else
		x"0000" when address_in = 16#00E9# else
		x"0000" when address_in = 16#00EA# else
		x"0000" when address_in = 16#00EB# else
		x"0000" when address_in = 16#00EC# else
		x"0000" when address_in = 16#00ED# else
		x"0000" when address_in = 16#00EE# else
		x"0000" when address_in = 16#00EF# else
		x"0000" when address_in = 16#00F0# else
		x"0000" when address_in = 16#00F1# else
		x"0000" when address_in = 16#00F2# else
		x"0000" when address_in = 16#00F3# else
		x"0000" when address_in = 16#00F4# else
		x"0000" when address_in = 16#00F5# else
		x"0000" when address_in = 16#00F6# else
		x"0000" when address_in = 16#00F7# else
		x"0000" when address_in = 16#00F8# else
		x"0000" when address_in = 16#00F9# else
		x"0000" when address_in = 16#00FA# else
		x"0000" when address_in = 16#00FB# else
		x"0000" when address_in = 16#00FC# else
		x"0000" when address_in = 16#00FD# else
		x"0000" when address_in = 16#00FE# else
		x"0000" when address_in = 16#00FF# else
		x"0000" when address_in = 16#0100# else
		x"0000" when address_in = 16#0101# else
		x"0000" when address_in = 16#0102# else
		x"0000" when address_in = 16#0103# else
		x"0000" when address_in = 16#0104# else
		x"0000" when address_in = 16#0105# else
		x"0000" when address_in = 16#0106# else
		x"0000" when address_in = 16#0107# else
		x"0000" when address_in = 16#0108# else
		x"0000" when address_in = 16#0109# else
		x"0000" when address_in = 16#010A# else
		x"0000" when address_in = 16#010B# else
		x"0000" when address_in = 16#010C# else
		x"0000" when address_in = 16#010D# else
		x"0000" when address_in = 16#010E# else
		x"0000" when address_in = 16#010F# else
		x"0000" when address_in = 16#0110# else
		x"0000" when address_in = 16#0111# else
		x"0000" when address_in = 16#0112# else
		x"0000" when address_in = 16#0113# else
		x"0000" when address_in = 16#0114# else
		x"0000" when address_in = 16#0115# else
		x"0000" when address_in = 16#0116# else
		x"0000" when address_in = 16#0117# else
		x"0000" when address_in = 16#0118# else
		x"0000" when address_in = 16#0119# else
		x"0000" when address_in = 16#011A# else
		x"0000" when address_in = 16#011B# else
		x"0000" when address_in = 16#011C# else
		x"0000" when address_in = 16#011D# else
		x"0000" when address_in = 16#011E# else
		x"0000" when address_in = 16#011F# else
		x"0000" when address_in = 16#0120# else
		x"0000" when address_in = 16#0121# else
		x"0000" when address_in = 16#0122# else
		x"0000" when address_in = 16#0123# else
		x"0000" when address_in = 16#0124# else
		x"0000" when address_in = 16#0125# else
		x"0000" when address_in = 16#0126# else
		x"0000" when address_in = 16#0127# else
		x"0000" when address_in = 16#0128# else
		x"0000" when address_in = 16#0129# else
		x"0000" when address_in = 16#012A# else
		x"0000" when address_in = 16#012B# else
		x"0000" when address_in = 16#012C# else
		x"0000" when address_in = 16#012D# else
		x"0000" when address_in = 16#012E# else
		x"0000" when address_in = 16#012F# else
		x"0000" when address_in = 16#0130# else
		x"0000" when address_in = 16#0131# else
		x"0000" when address_in = 16#0132# else
		x"0000" when address_in = 16#0133# else
		x"0000" when address_in = 16#0134# else
		x"0000" when address_in = 16#0135# else
		x"0000" when address_in = 16#0136# else
		x"0000" when address_in = 16#0137# else
		x"0000" when address_in = 16#0138# else
		x"0000" when address_in = 16#0139# else
		x"0000" when address_in = 16#013A# else
		x"0000" when address_in = 16#013B# else
		x"0000" when address_in = 16#013C# else
		x"0000" when address_in = 16#013D# else
		x"0000" when address_in = 16#013E# else
		x"0000" when address_in = 16#013F# else
		x"0000" when address_in = 16#0140# else
		x"0000" when address_in = 16#0141# else
		x"0000" when address_in = 16#0142# else
		x"0000" when address_in = 16#0143# else
		x"0000" when address_in = 16#0144# else
		x"0000" when address_in = 16#0145# else
		x"0000" when address_in = 16#0146# else
		x"0000" when address_in = 16#0147# else
		x"0000" when address_in = 16#0148# else
		x"0000" when address_in = 16#0149# else
		x"0000" when address_in = 16#014A# else
		x"0000" when address_in = 16#014B# else
		x"0000" when address_in = 16#014C# else
		x"0000" when address_in = 16#014D# else
		x"0000" when address_in = 16#014E# else
		x"0000" when address_in = 16#014F# else
		x"0000" when address_in = 16#0150# else
		x"0000" when address_in = 16#0151# else
		x"0000" when address_in = 16#0152# else
		x"0000" when address_in = 16#0153# else
		x"0000" when address_in = 16#0154# else
		x"0000" when address_in = 16#0155# else
		x"0000" when address_in = 16#0156# else
		x"0000" when address_in = 16#0157# else
		x"0000" when address_in = 16#0158# else
		x"0000" when address_in = 16#0159# else
		x"0000" when address_in = 16#015A# else
		x"0000" when address_in = 16#015B# else
		x"0000" when address_in = 16#015C# else
		x"0000" when address_in = 16#015D# else
		x"0000" when address_in = 16#015E# else
		x"0000" when address_in = 16#015F# else
		x"0000" when address_in = 16#0160# else
		x"0000" when address_in = 16#0161# else
		x"0000" when address_in = 16#0162# else
		x"0000" when address_in = 16#0163# else
		x"0000" when address_in = 16#0164# else
		x"0000" when address_in = 16#0165# else
		x"0000" when address_in = 16#0166# else
		x"0000" when address_in = 16#0167# else
		x"0000" when address_in = 16#0168# else
		x"0000" when address_in = 16#0169# else
		x"0000" when address_in = 16#016A# else
		x"0000" when address_in = 16#016B# else
		x"0000" when address_in = 16#016C# else
		x"0000" when address_in = 16#016D# else
		x"0000" when address_in = 16#016E# else
		x"0000" when address_in = 16#016F# else
		x"0000" when address_in = 16#0170# else
		x"0000" when address_in = 16#0171# else
		x"0000" when address_in = 16#0172# else
		x"0000" when address_in = 16#0173# else
		x"0000" when address_in = 16#0174# else
		x"0000" when address_in = 16#0175# else
		x"0000" when address_in = 16#0176# else
		x"0000" when address_in = 16#0177# else
		x"0000" when address_in = 16#0178# else
		x"0000" when address_in = 16#0179# else
		x"0000" when address_in = 16#017A# else
		x"0000" when address_in = 16#017B# else
		x"0000" when address_in = 16#017C# else
		x"0000" when address_in = 16#017D# else
		x"0000" when address_in = 16#017E# else
		x"0000" when address_in = 16#017F# else
		x"0000" when address_in = 16#0180# else
		x"0000" when address_in = 16#0181# else
		x"0000" when address_in = 16#0182# else
		x"0000" when address_in = 16#0183# else
		x"0000" when address_in = 16#0184# else
		x"0000" when address_in = 16#0185# else
		x"0000" when address_in = 16#0186# else
		x"0000" when address_in = 16#0187# else
		x"0000" when address_in = 16#0188# else
		x"0000" when address_in = 16#0189# else
		x"0000" when address_in = 16#018A# else
		x"0000" when address_in = 16#018B# else
		x"0000" when address_in = 16#018C# else
		x"0000" when address_in = 16#018D# else
		x"0000" when address_in = 16#018E# else
		x"0000" when address_in = 16#018F# else
		x"0000" when address_in = 16#0190# else
		x"0000" when address_in = 16#0191# else
		x"0000" when address_in = 16#0192# else
		x"0000" when address_in = 16#0193# else
		x"0000" when address_in = 16#0194# else
		x"0000" when address_in = 16#0195# else
		x"0000" when address_in = 16#0196# else
		x"0000" when address_in = 16#0197# else
		x"0000" when address_in = 16#0198# else
		x"0000" when address_in = 16#0199# else
		x"0000" when address_in = 16#019A# else
		x"0000" when address_in = 16#019B# else
		x"0000" when address_in = 16#019C# else
		x"0000" when address_in = 16#019D# else
		x"0000" when address_in = 16#019E# else
		x"0000" when address_in = 16#019F# else
		x"0000" when address_in = 16#01A0# else
		x"0000" when address_in = 16#01A1# else
		x"0000" when address_in = 16#01A2# else
		x"0000" when address_in = 16#01A3# else
		x"0000" when address_in = 16#01A4# else
		x"0000" when address_in = 16#01A5# else
		x"0000" when address_in = 16#01A6# else
		x"0000" when address_in = 16#01A7# else
		x"0000" when address_in = 16#01A8# else
		x"0000" when address_in = 16#01A9# else
		x"0000" when address_in = 16#01AA# else
		x"0000" when address_in = 16#01AB# else
		x"0000" when address_in = 16#01AC# else
		x"0000" when address_in = 16#01AD# else
		x"0000" when address_in = 16#01AE# else
		x"0000" when address_in = 16#01AF# else
		x"0000" when address_in = 16#01B0# else
		x"0000" when address_in = 16#01B1# else
		x"0000" when address_in = 16#01B2# else
		x"0000" when address_in = 16#01B3# else
		x"0000" when address_in = 16#01B4# else
		x"0000" when address_in = 16#01B5# else
		x"0000" when address_in = 16#01B6# else
		x"0000" when address_in = 16#01B7# else
		x"0000" when address_in = 16#01B8# else
		x"0000" when address_in = 16#01B9# else
		x"0000" when address_in = 16#01BA# else
		x"0000" when address_in = 16#01BB# else
		x"0000" when address_in = 16#01BC# else
		x"0000" when address_in = 16#01BD# else
		x"0000" when address_in = 16#01BE# else
		x"0000" when address_in = 16#01BF# else
		x"0000" when address_in = 16#01C0# else
		x"0000" when address_in = 16#01C1# else
		x"0000" when address_in = 16#01C2# else
		x"0000" when address_in = 16#01C3# else
		x"0000" when address_in = 16#01C4# else
		x"0000" when address_in = 16#01C5# else
		x"0000" when address_in = 16#01C6# else
		x"0000" when address_in = 16#01C7# else
		x"0000" when address_in = 16#01C8# else
		x"0000" when address_in = 16#01C9# else
		x"0000" when address_in = 16#01CA# else
		x"0000" when address_in = 16#01CB# else
		x"0000" when address_in = 16#01CC# else
		x"0000" when address_in = 16#01CD# else
		x"0000" when address_in = 16#01CE# else
		x"0000" when address_in = 16#01CF# else
		x"0000" when address_in = 16#01D0# else
		x"0000" when address_in = 16#01D1# else
		x"0000" when address_in = 16#01D2# else
		x"0000" when address_in = 16#01D3# else
		x"0000" when address_in = 16#01D4# else
		x"0000" when address_in = 16#01D5# else
		x"0000" when address_in = 16#01D6# else
		x"0000" when address_in = 16#01D7# else
		x"0000" when address_in = 16#01D8# else
		x"0000" when address_in = 16#01D9# else
		x"0000" when address_in = 16#01DA# else
		x"0000" when address_in = 16#01DB# else
		x"0000" when address_in = 16#01DC# else
		x"0000" when address_in = 16#01DD# else
		x"0000" when address_in = 16#01DE# else
		x"0000" when address_in = 16#01DF# else
		x"0000" when address_in = 16#01E0# else
		x"0000" when address_in = 16#01E1# else
		x"0000" when address_in = 16#01E2# else
		x"0000" when address_in = 16#01E3# else
		x"0000" when address_in = 16#01E4# else
		x"0000" when address_in = 16#01E5# else
		x"0000" when address_in = 16#01E6# else
		x"0000" when address_in = 16#01E7# else
		x"0000" when address_in = 16#01E8# else
		x"0000" when address_in = 16#01E9# else
		x"0000" when address_in = 16#01EA# else
		x"0000" when address_in = 16#01EB# else
		x"0000" when address_in = 16#01EC# else
		x"0000" when address_in = 16#01ED# else
		x"0000" when address_in = 16#01EE# else
		x"0000" when address_in = 16#01EF# else
		x"0000" when address_in = 16#01F0# else
		x"0000" when address_in = 16#01F1# else
		x"0000" when address_in = 16#01F2# else
		x"0000" when address_in = 16#01F3# else
		x"0000" when address_in = 16#01F4# else
		x"0000" when address_in = 16#01F5# else
		x"0000" when address_in = 16#01F6# else
		x"0000" when address_in = 16#01F7# else
		x"0000" when address_in = 16#01F8# else
		x"0000" when address_in = 16#01F9# else
		x"0000" when address_in = 16#01FA# else
		x"0000" when address_in = 16#01FB# else
		x"0000" when address_in = 16#01FC# else
		x"0000" when address_in = 16#01FD# else
		x"0000" when address_in = 16#01FE# else
		x"0000" when address_in = 16#01FF# else
		x"0000" when address_in = 16#0200# else
		x"0000" when address_in = 16#0201# else
		x"0000" when address_in = 16#0202# else
		x"0000" when address_in = 16#0203# else
		x"0000" when address_in = 16#0204# else
		x"0000" when address_in = 16#0205# else
		x"0000" when address_in = 16#0206# else
		x"0000" when address_in = 16#0207# else
		x"0000" when address_in = 16#0208# else
		x"0000" when address_in = 16#0209# else
		x"0000" when address_in = 16#020A# else
		x"0000" when address_in = 16#020B# else
		x"0000" when address_in = 16#020C# else
		x"0000" when address_in = 16#020D# else
		x"0000" when address_in = 16#020E# else
		x"0000" when address_in = 16#020F# else
		x"0000" when address_in = 16#0210# else
		x"0000" when address_in = 16#0211# else
		x"0000" when address_in = 16#0212# else
		x"0000" when address_in = 16#0213# else
		x"0000" when address_in = 16#0214# else
		x"0000" when address_in = 16#0215# else
		x"0000" when address_in = 16#0216# else
		x"0000" when address_in = 16#0217# else
		x"0000" when address_in = 16#0218# else
		x"0000" when address_in = 16#0219# else
		x"0000" when address_in = 16#021A# else
		x"0000" when address_in = 16#021B# else
		x"0000" when address_in = 16#021C# else
		x"0000" when address_in = 16#021D# else
		x"0000" when address_in = 16#021E# else
		x"0000" when address_in = 16#021F# else
		x"0000" when address_in = 16#0220# else
		x"0000" when address_in = 16#0221# else
		x"0000" when address_in = 16#0222# else
		x"0000" when address_in = 16#0223# else
		x"0000" when address_in = 16#0224# else
		x"0000" when address_in = 16#0225# else
		x"0000" when address_in = 16#0226# else
		x"0000" when address_in = 16#0227# else
		x"0000" when address_in = 16#0228# else
		x"0000" when address_in = 16#0229# else
		x"0000" when address_in = 16#022A# else
		x"0000" when address_in = 16#022B# else
		x"0000" when address_in = 16#022C# else
		x"0000" when address_in = 16#022D# else
		x"0000" when address_in = 16#022E# else
		x"0000" when address_in = 16#022F# else
		x"0000" when address_in = 16#0230# else
		x"0000" when address_in = 16#0231# else
		x"0000" when address_in = 16#0232# else
		x"0000" when address_in = 16#0233# else
		x"0000" when address_in = 16#0234# else
		x"0000" when address_in = 16#0235# else
		x"0000" when address_in = 16#0236# else
		x"0000" when address_in = 16#0237# else
		x"0000" when address_in = 16#0238# else
		x"0000" when address_in = 16#0239# else
		x"0000" when address_in = 16#023A# else
		x"0000" when address_in = 16#023B# else
		x"0000" when address_in = 16#023C# else
		x"0000" when address_in = 16#023D# else
		x"0000" when address_in = 16#023E# else
		x"0000" when address_in = 16#023F# else
		x"0000" when address_in = 16#0240# else
		x"0000" when address_in = 16#0241# else
		x"0000" when address_in = 16#0242# else
		x"0000" when address_in = 16#0243# else
		x"0000" when address_in = 16#0244# else
		x"0000" when address_in = 16#0245# else
		x"0000" when address_in = 16#0246# else
		x"0000" when address_in = 16#0247# else
		x"0000" when address_in = 16#0248# else
		x"0000" when address_in = 16#0249# else
		x"0000" when address_in = 16#024A# else
		x"0000" when address_in = 16#024B# else
		x"0000" when address_in = 16#024C# else
		x"0000" when address_in = 16#024D# else
		x"0000" when address_in = 16#024E# else
		x"0000" when address_in = 16#024F# else
		x"0000" when address_in = 16#0250# else
		x"0000" when address_in = 16#0251# else
		x"0000" when address_in = 16#0252# else
		x"0000" when address_in = 16#0253# else
		x"0000" when address_in = 16#0254# else
		x"0000" when address_in = 16#0255# else
		x"0000" when address_in = 16#0256# else
		x"0000" when address_in = 16#0257# else
		x"0000" when address_in = 16#0258# else
		x"0000" when address_in = 16#0259# else
		x"0000" when address_in = 16#025A# else
		x"0000" when address_in = 16#025B# else
		x"0000" when address_in = 16#025C# else
		x"0000" when address_in = 16#025D# else
		x"0000" when address_in = 16#025E# else
		x"0000" when address_in = 16#025F# else
		x"0000" when address_in = 16#0260# else
		x"0000" when address_in = 16#0261# else
		x"0000" when address_in = 16#0262# else
		x"0000" when address_in = 16#0263# else
		x"0000" when address_in = 16#0264# else
		x"0000" when address_in = 16#0265# else
		x"0000" when address_in = 16#0266# else
		x"0000" when address_in = 16#0267# else
		x"0000" when address_in = 16#0268# else
		x"0000" when address_in = 16#0269# else
		x"0000" when address_in = 16#026A# else
		x"0000" when address_in = 16#026B# else
		x"0000" when address_in = 16#026C# else
		x"0000" when address_in = 16#026D# else
		x"0000" when address_in = 16#026E# else
		x"0000" when address_in = 16#026F# else
		x"0000" when address_in = 16#0270# else
		x"0000" when address_in = 16#0271# else
		x"0000" when address_in = 16#0272# else
		x"0000" when address_in = 16#0273# else
		x"0000" when address_in = 16#0274# else
		x"0000" when address_in = 16#0275# else
		x"0000" when address_in = 16#0276# else
		x"0000" when address_in = 16#0277# else
		x"0000" when address_in = 16#0278# else
		x"0000" when address_in = 16#0279# else
		x"0000" when address_in = 16#027A# else
		x"0000" when address_in = 16#027B# else
		x"0000" when address_in = 16#027C# else
		x"0000" when address_in = 16#027D# else
		x"0000" when address_in = 16#027E# else
		x"0000" when address_in = 16#027F# else
		x"0000" when address_in = 16#0280# else
		x"0000" when address_in = 16#0281# else
		x"0000" when address_in = 16#0282# else
		x"0000" when address_in = 16#0283# else
		x"0000" when address_in = 16#0284# else
		x"0000" when address_in = 16#0285# else
		x"0000" when address_in = 16#0286# else
		x"0000" when address_in = 16#0287# else
		x"0000" when address_in = 16#0288# else
		x"0000" when address_in = 16#0289# else
		x"0000" when address_in = 16#028A# else
		x"0000" when address_in = 16#028B# else
		x"0000" when address_in = 16#028C# else
		x"0000" when address_in = 16#028D# else
		x"0000" when address_in = 16#028E# else
		x"0000" when address_in = 16#028F# else
		x"0000" when address_in = 16#0290# else
		x"0000" when address_in = 16#0291# else
		x"0000" when address_in = 16#0292# else
		x"0000" when address_in = 16#0293# else
		x"0000" when address_in = 16#0294# else
		x"0000" when address_in = 16#0295# else
		x"0000" when address_in = 16#0296# else
		x"0000" when address_in = 16#0297# else
		x"0000" when address_in = 16#0298# else
		x"0000" when address_in = 16#0299# else
		x"0000" when address_in = 16#029A# else
		x"0000" when address_in = 16#029B# else
		x"0000" when address_in = 16#029C# else
		x"0000" when address_in = 16#029D# else
		x"0000" when address_in = 16#029E# else
		x"0000" when address_in = 16#029F# else
		x"0000" when address_in = 16#02A0# else
		x"0000" when address_in = 16#02A1# else
		x"0000" when address_in = 16#02A2# else
		x"0000" when address_in = 16#02A3# else
		x"0000" when address_in = 16#02A4# else
		x"0000" when address_in = 16#02A5# else
		x"0000" when address_in = 16#02A6# else
		x"0000" when address_in = 16#02A7# else
		x"0000" when address_in = 16#02A8# else
		x"0000" when address_in = 16#02A9# else
		x"0000" when address_in = 16#02AA# else
		x"0000" when address_in = 16#02AB# else
		x"0000" when address_in = 16#02AC# else
		x"0000" when address_in = 16#02AD# else
		x"0000" when address_in = 16#02AE# else
		x"0000" when address_in = 16#02AF# else
		x"0000" when address_in = 16#02B0# else
		x"0000" when address_in = 16#02B1# else
		x"0000" when address_in = 16#02B2# else
		x"0000" when address_in = 16#02B3# else
		x"0000" when address_in = 16#02B4# else
		x"0000" when address_in = 16#02B5# else
		x"0000" when address_in = 16#02B6# else
		x"0000" when address_in = 16#02B7# else
		x"0000" when address_in = 16#02B8# else
		x"0000" when address_in = 16#02B9# else
		x"0000" when address_in = 16#02BA# else
		x"0000" when address_in = 16#02BB# else
		x"0000" when address_in = 16#02BC# else
		x"0000" when address_in = 16#02BD# else
		x"0000" when address_in = 16#02BE# else
		x"0000" when address_in = 16#02BF# else
		x"0000" when address_in = 16#02C0# else
		x"0000" when address_in = 16#02C1# else
		x"0000" when address_in = 16#02C2# else
		x"0000" when address_in = 16#02C3# else
		x"0000" when address_in = 16#02C4# else
		x"0000" when address_in = 16#02C5# else
		x"0000" when address_in = 16#02C6# else
		x"0000" when address_in = 16#02C7# else
		x"0000" when address_in = 16#02C8# else
		x"0000" when address_in = 16#02C9# else
		x"0000" when address_in = 16#02CA# else
		x"0000" when address_in = 16#02CB# else
		x"0000" when address_in = 16#02CC# else
		x"0000" when address_in = 16#02CD# else
		x"0000" when address_in = 16#02CE# else
		x"0000" when address_in = 16#02CF# else
		x"0000" when address_in = 16#02D0# else
		x"0000" when address_in = 16#02D1# else
		x"0000" when address_in = 16#02D2# else
		x"0000" when address_in = 16#02D3# else
		x"0000" when address_in = 16#02D4# else
		x"0000" when address_in = 16#02D5# else
		x"0000" when address_in = 16#02D6# else
		x"0000" when address_in = 16#02D7# else
		x"0000" when address_in = 16#02D8# else
		x"0000" when address_in = 16#02D9# else
		x"0000" when address_in = 16#02DA# else
		x"0000" when address_in = 16#02DB# else
		x"0000" when address_in = 16#02DC# else
		x"0000" when address_in = 16#02DD# else
		x"0000" when address_in = 16#02DE# else
		x"0000" when address_in = 16#02DF# else
		x"0000" when address_in = 16#02E0# else
		x"0000" when address_in = 16#02E1# else
		x"0000" when address_in = 16#02E2# else
		x"0000" when address_in = 16#02E3# else
		x"0000" when address_in = 16#02E4# else
		x"0000" when address_in = 16#02E5# else
		x"0000" when address_in = 16#02E6# else
		x"0000" when address_in = 16#02E7# else
		x"0000" when address_in = 16#02E8# else
		x"0000" when address_in = 16#02E9# else
		x"0000" when address_in = 16#02EA# else
		x"0000" when address_in = 16#02EB# else
		x"0000" when address_in = 16#02EC# else
		x"0000" when address_in = 16#02ED# else
		x"0000" when address_in = 16#02EE# else
		x"0000" when address_in = 16#02EF# else
		x"0000" when address_in = 16#02F0# else
		x"0000" when address_in = 16#02F1# else
		x"0000" when address_in = 16#02F2# else
		x"0000" when address_in = 16#02F3# else
		x"0000" when address_in = 16#02F4# else
		x"0000" when address_in = 16#02F5# else
		x"0000" when address_in = 16#02F6# else
		x"0000" when address_in = 16#02F7# else
		x"0000" when address_in = 16#02F8# else
		x"0000" when address_in = 16#02F9# else
		x"0000" when address_in = 16#02FA# else
		x"0000" when address_in = 16#02FB# else
		x"0000" when address_in = 16#02FC# else
		x"0000" when address_in = 16#02FD# else
		x"0000" when address_in = 16#02FE# else
		x"0000" when address_in = 16#02FF# else
		x"0000" when address_in = 16#0300# else
		x"0000" when address_in = 16#0301# else
		x"0000" when address_in = 16#0302# else
		x"0000" when address_in = 16#0303# else
		x"0000" when address_in = 16#0304# else
		x"0000" when address_in = 16#0305# else
		x"0000" when address_in = 16#0306# else
		x"0000" when address_in = 16#0307# else
		x"0000" when address_in = 16#0308# else
		x"0000" when address_in = 16#0309# else
		x"0000" when address_in = 16#030A# else
		x"0000" when address_in = 16#030B# else
		x"0000" when address_in = 16#030C# else
		x"0000" when address_in = 16#030D# else
		x"0000" when address_in = 16#030E# else
		x"0000" when address_in = 16#030F# else
		x"0000" when address_in = 16#0310# else
		x"0000" when address_in = 16#0311# else
		x"0000" when address_in = 16#0312# else
		x"0000" when address_in = 16#0313# else
		x"0000" when address_in = 16#0314# else
		x"0000" when address_in = 16#0315# else
		x"0000" when address_in = 16#0316# else
		x"0000" when address_in = 16#0317# else
		x"0000" when address_in = 16#0318# else
		x"0000" when address_in = 16#0319# else
		x"0000" when address_in = 16#031A# else
		x"0000" when address_in = 16#031B# else
		x"0000" when address_in = 16#031C# else
		x"0000" when address_in = 16#031D# else
		x"0000" when address_in = 16#031E# else
		x"0000" when address_in = 16#031F# else
		x"0000" when address_in = 16#0320# else
		x"0000" when address_in = 16#0321# else
		x"0000" when address_in = 16#0322# else
		x"0000" when address_in = 16#0323# else
		x"0000" when address_in = 16#0324# else
		x"0000" when address_in = 16#0325# else
		x"0000" when address_in = 16#0326# else
		x"0000" when address_in = 16#0327# else
		x"0000" when address_in = 16#0328# else
		x"0000" when address_in = 16#0329# else
		x"0000" when address_in = 16#032A# else
		x"0000" when address_in = 16#032B# else
		x"0000" when address_in = 16#032C# else
		x"0000" when address_in = 16#032D# else
		x"0000" when address_in = 16#032E# else
		x"0000" when address_in = 16#032F# else
		x"0000" when address_in = 16#0330# else
		x"0000" when address_in = 16#0331# else
		x"0000" when address_in = 16#0332# else
		x"0000" when address_in = 16#0333# else
		x"0000" when address_in = 16#0334# else
		x"0000" when address_in = 16#0335# else
		x"0000" when address_in = 16#0336# else
		x"0000" when address_in = 16#0337# else
		x"0000" when address_in = 16#0338# else
		x"0000" when address_in = 16#0339# else
		x"0000" when address_in = 16#033A# else
		x"0000" when address_in = 16#033B# else
		x"0000" when address_in = 16#033C# else
		x"0000" when address_in = 16#033D# else
		x"0000" when address_in = 16#033E# else
		x"0000" when address_in = 16#033F# else
		x"0000" when address_in = 16#0340# else
		x"0000" when address_in = 16#0341# else
		x"0000" when address_in = 16#0342# else
		x"0000" when address_in = 16#0343# else
		x"0000" when address_in = 16#0344# else
		x"0000" when address_in = 16#0345# else
		x"0000" when address_in = 16#0346# else
		x"0000" when address_in = 16#0347# else
		x"0000" when address_in = 16#0348# else
		x"0000" when address_in = 16#0349# else
		x"0000" when address_in = 16#034A# else
		x"0000" when address_in = 16#034B# else
		x"0000" when address_in = 16#034C# else
		x"0000" when address_in = 16#034D# else
		x"0000" when address_in = 16#034E# else
		x"0000" when address_in = 16#034F# else
		x"0000" when address_in = 16#0350# else
		x"0000" when address_in = 16#0351# else
		x"0000" when address_in = 16#0352# else
		x"0000" when address_in = 16#0353# else
		x"0000" when address_in = 16#0354# else
		x"0000" when address_in = 16#0355# else
		x"0000" when address_in = 16#0356# else
		x"0000" when address_in = 16#0357# else
		x"0000" when address_in = 16#0358# else
		x"0000" when address_in = 16#0359# else
		x"0000" when address_in = 16#035A# else
		x"0000" when address_in = 16#035B# else
		x"0000" when address_in = 16#035C# else
		x"0000" when address_in = 16#035D# else
		x"0000" when address_in = 16#035E# else
		x"0000" when address_in = 16#035F# else
		x"0000" when address_in = 16#0360# else
		x"0000" when address_in = 16#0361# else
		x"0000" when address_in = 16#0362# else
		x"0000" when address_in = 16#0363# else
		x"0000" when address_in = 16#0364# else
		x"0000" when address_in = 16#0365# else
		x"0000" when address_in = 16#0366# else
		x"0000" when address_in = 16#0367# else
		x"0000" when address_in = 16#0368# else
		x"0000" when address_in = 16#0369# else
		x"0000" when address_in = 16#036A# else
		x"0000" when address_in = 16#036B# else
		x"0000" when address_in = 16#036C# else
		x"0000" when address_in = 16#036D# else
		x"0000" when address_in = 16#036E# else
		x"0000" when address_in = 16#036F# else
		x"0000" when address_in = 16#0370# else
		x"0000" when address_in = 16#0371# else
		x"0000" when address_in = 16#0372# else
		x"0000" when address_in = 16#0373# else
		x"0000" when address_in = 16#0374# else
		x"0000" when address_in = 16#0375# else
		x"0000" when address_in = 16#0376# else
		x"0000" when address_in = 16#0377# else
		x"0000" when address_in = 16#0378# else
		x"0000" when address_in = 16#0379# else
		x"0000" when address_in = 16#037A# else
		x"0000" when address_in = 16#037B# else
		x"0000" when address_in = 16#037C# else
		x"0000" when address_in = 16#037D# else
		x"0000" when address_in = 16#037E# else
		x"0000" when address_in = 16#037F# else
		x"0000" when address_in = 16#0380# else
		x"0000" when address_in = 16#0381# else
		x"0000" when address_in = 16#0382# else
		x"0000" when address_in = 16#0383# else
		x"0000" when address_in = 16#0384# else
		x"0000" when address_in = 16#0385# else
		x"0000" when address_in = 16#0386# else
		x"0000" when address_in = 16#0387# else
		x"0000" when address_in = 16#0388# else
		x"0000" when address_in = 16#0389# else
		x"0000" when address_in = 16#038A# else
		x"0000" when address_in = 16#038B# else
		x"0000" when address_in = 16#038C# else
		x"0000" when address_in = 16#038D# else
		x"0000" when address_in = 16#038E# else
		x"0000" when address_in = 16#038F# else
		x"0000" when address_in = 16#0390# else
		x"0000" when address_in = 16#0391# else
		x"0000" when address_in = 16#0392# else
		x"0000" when address_in = 16#0393# else
		x"0000" when address_in = 16#0394# else
		x"0000" when address_in = 16#0395# else
		x"0000" when address_in = 16#0396# else
		x"0000" when address_in = 16#0397# else
		x"0000" when address_in = 16#0398# else
		x"0000" when address_in = 16#0399# else
		x"0000" when address_in = 16#039A# else
		x"0000" when address_in = 16#039B# else
		x"0000" when address_in = 16#039C# else
		x"0000" when address_in = 16#039D# else
		x"0000" when address_in = 16#039E# else
		x"0000" when address_in = 16#039F# else
		x"0000" when address_in = 16#03A0# else
		x"0000" when address_in = 16#03A1# else
		x"0000" when address_in = 16#03A2# else
		x"0000" when address_in = 16#03A3# else
		x"0000" when address_in = 16#03A4# else
		x"0000" when address_in = 16#03A5# else
		x"0000" when address_in = 16#03A6# else
		x"0000" when address_in = 16#03A7# else
		x"0000" when address_in = 16#03A8# else
		x"0000" when address_in = 16#03A9# else
		x"0000" when address_in = 16#03AA# else
		x"0000" when address_in = 16#03AB# else
		x"0000" when address_in = 16#03AC# else
		x"0000" when address_in = 16#03AD# else
		x"0000" when address_in = 16#03AE# else
		x"0000" when address_in = 16#03AF# else
		x"0000" when address_in = 16#03B0# else
		x"0000" when address_in = 16#03B1# else
		x"0000" when address_in = 16#03B2# else
		x"0000" when address_in = 16#03B3# else
		x"0000" when address_in = 16#03B4# else
		x"0000" when address_in = 16#03B5# else
		x"0000" when address_in = 16#03B6# else
		x"0000" when address_in = 16#03B7# else
		x"0000" when address_in = 16#03B8# else
		x"0000" when address_in = 16#03B9# else
		x"0000" when address_in = 16#03BA# else
		x"0000" when address_in = 16#03BB# else
		x"0000" when address_in = 16#03BC# else
		x"0000" when address_in = 16#03BD# else
		x"0000" when address_in = 16#03BE# else
		x"0000" when address_in = 16#03BF# else
		x"0000" when address_in = 16#03C0# else
		x"0000" when address_in = 16#03C1# else
		x"0000" when address_in = 16#03C2# else
		x"0000" when address_in = 16#03C3# else
		x"0000" when address_in = 16#03C4# else
		x"0000" when address_in = 16#03C5# else
		x"0000" when address_in = 16#03C6# else
		x"0000" when address_in = 16#03C7# else
		x"0000" when address_in = 16#03C8# else
		x"0000" when address_in = 16#03C9# else
		x"0000" when address_in = 16#03CA# else
		x"0000" when address_in = 16#03CB# else
		x"0000" when address_in = 16#03CC# else
		x"0000" when address_in = 16#03CD# else
		x"0000" when address_in = 16#03CE# else
		x"0000" when address_in = 16#03CF# else
		x"0000" when address_in = 16#03D0# else
		x"0000" when address_in = 16#03D1# else
		x"0000" when address_in = 16#03D2# else
		x"0000" when address_in = 16#03D3# else
		x"0000" when address_in = 16#03D4# else
		x"0000" when address_in = 16#03D5# else
		x"0000" when address_in = 16#03D6# else
		x"0000" when address_in = 16#03D7# else
		x"0000" when address_in = 16#03D8# else
		x"0000" when address_in = 16#03D9# else
		x"0000" when address_in = 16#03DA# else
		x"0000" when address_in = 16#03DB# else
		x"0000" when address_in = 16#03DC# else
		x"0000" when address_in = 16#03DD# else
		x"0000" when address_in = 16#03DE# else
		x"0000" when address_in = 16#03DF# else
		x"0000" when address_in = 16#03E0# else
		x"0000" when address_in = 16#03E1# else
		x"0000" when address_in = 16#03E2# else
		x"0000" when address_in = 16#03E3# else
		x"0000" when address_in = 16#03E4# else
		x"0000" when address_in = 16#03E5# else
		x"0000" when address_in = 16#03E6# else
		x"0000" when address_in = 16#03E7# else
		x"0000" when address_in = 16#03E8# else
		x"0000" when address_in = 16#03E9# else
		x"0000" when address_in = 16#03EA# else
		x"0000" when address_in = 16#03EB# else
		x"0000" when address_in = 16#03EC# else
		x"0000" when address_in = 16#03ED# else
		x"0000" when address_in = 16#03EE# else
		x"0000" when address_in = 16#03EF# else
		x"0000" when address_in = 16#03F0# else
		x"0000" when address_in = 16#03F1# else
		x"0000" when address_in = 16#03F2# else
		x"0000" when address_in = 16#03F3# else
		x"0000" when address_in = 16#03F4# else
		x"0000" when address_in = 16#03F5# else
		x"0000" when address_in = 16#03F6# else
		x"0000" when address_in = 16#03F7# else
		x"0000" when address_in = 16#03F8# else
		x"0000" when address_in = 16#03F9# else
		x"0000" when address_in = 16#03FA# else
		x"0000" when address_in = 16#03FB# else
		x"0000" when address_in = 16#03FC# else
		x"0000" when address_in = 16#03FD# else
		x"0000" when address_in = 16#03FE# else
		x"0000" when address_in = 16#03FF# else
		x"940C" when address_in = 16#0400# else
		x"2E2C" when address_in = 16#0401# else
		x"940C" when address_in = 16#0402# else
		x"0A00" when address_in = 16#0403# else
		x"940C" when address_in = 16#0404# else
		x"0000" when address_in = 16#0405# else
		x"940C" when address_in = 16#0406# else
		x"0A22" when address_in = 16#0407# else
		x"940C" when address_in = 16#0408# else
		x"10FC" when address_in = 16#0409# else
		x"940C" when address_in = 16#040A# else
		x"2027" when address_in = 16#040B# else
		x"940C" when address_in = 16#040C# else
		x"2058" when address_in = 16#040D# else
		x"940C" when address_in = 16#040E# else
		x"207F" when address_in = 16#040F# else
		x"940C" when address_in = 16#0410# else
		x"1078" when address_in = 16#0411# else
		x"940C" when address_in = 16#0412# else
		x"1503" when address_in = 16#0413# else
		x"940C" when address_in = 16#0414# else
		x"1119" when address_in = 16#0415# else
		x"940C" when address_in = 16#0416# else
		x"255D" when address_in = 16#0417# else
		x"940C" when address_in = 16#0418# else
		x"2433" when address_in = 16#0419# else
		x"940C" when address_in = 16#041A# else
		x"258C" when address_in = 16#041B# else
		x"940C" when address_in = 16#041C# else
		x"0000" when address_in = 16#041D# else
		x"940C" when address_in = 16#041E# else
		x"0000" when address_in = 16#041F# else
		x"940C" when address_in = 16#0420# else
		x"26CF" when address_in = 16#0421# else
		x"940C" when address_in = 16#0422# else
		x"0B48" when address_in = 16#0423# else
		x"940C" when address_in = 16#0424# else
		x"1B46" when address_in = 16#0425# else
		x"940C" when address_in = 16#0426# else
		x"0A25" when address_in = 16#0427# else
		x"940C" when address_in = 16#0428# else
		x"0000" when address_in = 16#0429# else
		x"940C" when address_in = 16#042A# else
		x"0000" when address_in = 16#042B# else
		x"940C" when address_in = 16#042C# else
		x"0000" when address_in = 16#042D# else
		x"940C" when address_in = 16#042E# else
		x"0000" when address_in = 16#042F# else
		x"940C" when address_in = 16#0430# else
		x"0000" when address_in = 16#0431# else
		x"940C" when address_in = 16#0432# else
		x"0000" when address_in = 16#0433# else
		x"940C" when address_in = 16#0434# else
		x"0000" when address_in = 16#0435# else
		x"940C" when address_in = 16#0436# else
		x"0000" when address_in = 16#0437# else
		x"940C" when address_in = 16#0438# else
		x"0000" when address_in = 16#0439# else
		x"940C" when address_in = 16#043A# else
		x"0000" when address_in = 16#043B# else
		x"940C" when address_in = 16#043C# else
		x"0000" when address_in = 16#043D# else
		x"940C" when address_in = 16#043E# else
		x"0000" when address_in = 16#043F# else
		x"0000" when address_in = 16#0440# else
		x"0000" when address_in = 16#0441# else
		x"0000" when address_in = 16#0442# else
		x"0000" when address_in = 16#0443# else
		x"0000" when address_in = 16#0444# else
		x"0000" when address_in = 16#0445# else
		x"0000" when address_in = 16#0446# else
		x"0000" when address_in = 16#0447# else
		x"0000" when address_in = 16#0448# else
		x"0000" when address_in = 16#0449# else
		x"0000" when address_in = 16#044A# else
		x"0000" when address_in = 16#044B# else
		x"0000" when address_in = 16#044C# else
		x"0000" when address_in = 16#044D# else
		x"0000" when address_in = 16#044E# else
		x"0000" when address_in = 16#044F# else
		x"0000" when address_in = 16#0450# else
		x"0000" when address_in = 16#0451# else
		x"0000" when address_in = 16#0452# else
		x"0000" when address_in = 16#0453# else
		x"0000" when address_in = 16#0454# else
		x"0000" when address_in = 16#0455# else
		x"0000" when address_in = 16#0456# else
		x"0000" when address_in = 16#0457# else
		x"0000" when address_in = 16#0458# else
		x"0000" when address_in = 16#0459# else
		x"0000" when address_in = 16#045A# else
		x"0000" when address_in = 16#045B# else
		x"0000" when address_in = 16#045C# else
		x"0000" when address_in = 16#045D# else
		x"0000" when address_in = 16#045E# else
		x"0000" when address_in = 16#045F# else
		x"0000" when address_in = 16#0460# else
		x"0000" when address_in = 16#0461# else
		x"0000" when address_in = 16#0462# else
		x"0000" when address_in = 16#0463# else
		x"0000" when address_in = 16#0464# else
		x"0000" when address_in = 16#0465# else
		x"0000" when address_in = 16#0466# else
		x"0000" when address_in = 16#0467# else
		x"0000" when address_in = 16#0468# else
		x"0000" when address_in = 16#0469# else
		x"0000" when address_in = 16#046A# else
		x"0000" when address_in = 16#046B# else
		x"0000" when address_in = 16#046C# else
		x"0000" when address_in = 16#046D# else
		x"0000" when address_in = 16#046E# else
		x"0000" when address_in = 16#046F# else
		x"0000" when address_in = 16#0470# else
		x"0000" when address_in = 16#0471# else
		x"0000" when address_in = 16#0472# else
		x"0000" when address_in = 16#0473# else
		x"0000" when address_in = 16#0474# else
		x"0000" when address_in = 16#0475# else
		x"0000" when address_in = 16#0476# else
		x"0000" when address_in = 16#0477# else
		x"0000" when address_in = 16#0478# else
		x"0000" when address_in = 16#0479# else
		x"0000" when address_in = 16#047A# else
		x"0000" when address_in = 16#047B# else
		x"0000" when address_in = 16#047C# else
		x"0000" when address_in = 16#047D# else
		x"0000" when address_in = 16#047E# else
		x"0000" when address_in = 16#047F# else
		x"0280" when address_in = 16#0480# else
		x"0000" when address_in = 16#0481# else
		x"0000" when address_in = 16#0482# else
		x"0101" when address_in = 16#0483# else
		x"0080" when address_in = 16#0484# else
		x"0000" when address_in = 16#0485# else
		x"0080" when address_in = 16#0486# else
		x"0002" when address_in = 16#0487# else
		x"0000" when address_in = 16#0488# else
		x"0000" when address_in = 16#0489# else
		x"0000" when address_in = 16#048A# else
		x"0000" when address_in = 16#048B# else
		x"0007" when address_in = 16#048C# else
		x"0B0F" when address_in = 16#048D# else
		x"0048" when address_in = 16#048E# else
		x"0001" when address_in = 16#048F# else
		x"0000" when address_in = 16#0490# else
		x"0000" when address_in = 16#0491# else
		x"0000" when address_in = 16#0492# else
		x"0007" when address_in = 16#0493# else
		x"2629" when address_in = 16#0494# else
		x"0000" when address_in = 16#0495# else
		x"1021" when address_in = 16#0496# else
		x"2042" when address_in = 16#0497# else
		x"3063" when address_in = 16#0498# else
		x"4084" when address_in = 16#0499# else
		x"50A5" when address_in = 16#049A# else
		x"60C6" when address_in = 16#049B# else
		x"70E7" when address_in = 16#049C# else
		x"8108" when address_in = 16#049D# else
		x"9129" when address_in = 16#049E# else
		x"A14A" when address_in = 16#049F# else
		x"B16B" when address_in = 16#04A0# else
		x"C18C" when address_in = 16#04A1# else
		x"D1AD" when address_in = 16#04A2# else
		x"E1CE" when address_in = 16#04A3# else
		x"F1EF" when address_in = 16#04A4# else
		x"1231" when address_in = 16#04A5# else
		x"0210" when address_in = 16#04A6# else
		x"3273" when address_in = 16#04A7# else
		x"2252" when address_in = 16#04A8# else
		x"52B5" when address_in = 16#04A9# else
		x"4294" when address_in = 16#04AA# else
		x"72F7" when address_in = 16#04AB# else
		x"62D6" when address_in = 16#04AC# else
		x"9339" when address_in = 16#04AD# else
		x"8318" when address_in = 16#04AE# else
		x"B37B" when address_in = 16#04AF# else
		x"A35A" when address_in = 16#04B0# else
		x"D3BD" when address_in = 16#04B1# else
		x"C39C" when address_in = 16#04B2# else
		x"F3FF" when address_in = 16#04B3# else
		x"E3DE" when address_in = 16#04B4# else
		x"2462" when address_in = 16#04B5# else
		x"3443" when address_in = 16#04B6# else
		x"0420" when address_in = 16#04B7# else
		x"1401" when address_in = 16#04B8# else
		x"64E6" when address_in = 16#04B9# else
		x"74C7" when address_in = 16#04BA# else
		x"44A4" when address_in = 16#04BB# else
		x"5485" when address_in = 16#04BC# else
		x"A56A" when address_in = 16#04BD# else
		x"B54B" when address_in = 16#04BE# else
		x"8528" when address_in = 16#04BF# else
		x"9509" when address_in = 16#04C0# else
		x"E5EE" when address_in = 16#04C1# else
		x"F5CF" when address_in = 16#04C2# else
		x"C5AC" when address_in = 16#04C3# else
		x"D58D" when address_in = 16#04C4# else
		x"3653" when address_in = 16#04C5# else
		x"2672" when address_in = 16#04C6# else
		x"1611" when address_in = 16#04C7# else
		x"0630" when address_in = 16#04C8# else
		x"76D7" when address_in = 16#04C9# else
		x"66F6" when address_in = 16#04CA# else
		x"5695" when address_in = 16#04CB# else
		x"46B4" when address_in = 16#04CC# else
		x"B75B" when address_in = 16#04CD# else
		x"A77A" when address_in = 16#04CE# else
		x"9719" when address_in = 16#04CF# else
		x"8738" when address_in = 16#04D0# else
		x"F7DF" when address_in = 16#04D1# else
		x"E7FE" when address_in = 16#04D2# else
		x"D79D" when address_in = 16#04D3# else
		x"C7BC" when address_in = 16#04D4# else
		x"48C4" when address_in = 16#04D5# else
		x"58E5" when address_in = 16#04D6# else
		x"6886" when address_in = 16#04D7# else
		x"78A7" when address_in = 16#04D8# else
		x"0840" when address_in = 16#04D9# else
		x"1861" when address_in = 16#04DA# else
		x"2802" when address_in = 16#04DB# else
		x"3823" when address_in = 16#04DC# else
		x"C9CC" when address_in = 16#04DD# else
		x"D9ED" when address_in = 16#04DE# else
		x"E98E" when address_in = 16#04DF# else
		x"F9AF" when address_in = 16#04E0# else
		x"8948" when address_in = 16#04E1# else
		x"9969" when address_in = 16#04E2# else
		x"A90A" when address_in = 16#04E3# else
		x"B92B" when address_in = 16#04E4# else
		x"5AF5" when address_in = 16#04E5# else
		x"4AD4" when address_in = 16#04E6# else
		x"7AB7" when address_in = 16#04E7# else
		x"6A96" when address_in = 16#04E8# else
		x"1A71" when address_in = 16#04E9# else
		x"0A50" when address_in = 16#04EA# else
		x"3A33" when address_in = 16#04EB# else
		x"2A12" when address_in = 16#04EC# else
		x"DBFD" when address_in = 16#04ED# else
		x"CBDC" when address_in = 16#04EE# else
		x"FBBF" when address_in = 16#04EF# else
		x"EB9E" when address_in = 16#04F0# else
		x"9B79" when address_in = 16#04F1# else
		x"8B58" when address_in = 16#04F2# else
		x"BB3B" when address_in = 16#04F3# else
		x"AB1A" when address_in = 16#04F4# else
		x"6CA6" when address_in = 16#04F5# else
		x"7C87" when address_in = 16#04F6# else
		x"4CE4" when address_in = 16#04F7# else
		x"5CC5" when address_in = 16#04F8# else
		x"2C22" when address_in = 16#04F9# else
		x"3C03" when address_in = 16#04FA# else
		x"0C60" when address_in = 16#04FB# else
		x"1C41" when address_in = 16#04FC# else
		x"EDAE" when address_in = 16#04FD# else
		x"FD8F" when address_in = 16#04FE# else
		x"CDEC" when address_in = 16#04FF# else
		x"DDCD" when address_in = 16#0500# else
		x"AD2A" when address_in = 16#0501# else
		x"BD0B" when address_in = 16#0502# else
		x"8D68" when address_in = 16#0503# else
		x"9D49" when address_in = 16#0504# else
		x"7E97" when address_in = 16#0505# else
		x"6EB6" when address_in = 16#0506# else
		x"5ED5" when address_in = 16#0507# else
		x"4EF4" when address_in = 16#0508# else
		x"3E13" when address_in = 16#0509# else
		x"2E32" when address_in = 16#050A# else
		x"1E51" when address_in = 16#050B# else
		x"0E70" when address_in = 16#050C# else
		x"FF9F" when address_in = 16#050D# else
		x"EFBE" when address_in = 16#050E# else
		x"DFDD" when address_in = 16#050F# else
		x"CFFC" when address_in = 16#0510# else
		x"BF1B" when address_in = 16#0511# else
		x"AF3A" when address_in = 16#0512# else
		x"9F59" when address_in = 16#0513# else
		x"8F78" when address_in = 16#0514# else
		x"9188" when address_in = 16#0515# else
		x"81A9" when address_in = 16#0516# else
		x"B1CA" when address_in = 16#0517# else
		x"A1EB" when address_in = 16#0518# else
		x"D10C" when address_in = 16#0519# else
		x"C12D" when address_in = 16#051A# else
		x"F14E" when address_in = 16#051B# else
		x"E16F" when address_in = 16#051C# else
		x"1080" when address_in = 16#051D# else
		x"00A1" when address_in = 16#051E# else
		x"30C2" when address_in = 16#051F# else
		x"20E3" when address_in = 16#0520# else
		x"5004" when address_in = 16#0521# else
		x"4025" when address_in = 16#0522# else
		x"7046" when address_in = 16#0523# else
		x"6067" when address_in = 16#0524# else
		x"83B9" when address_in = 16#0525# else
		x"9398" when address_in = 16#0526# else
		x"A3FB" when address_in = 16#0527# else
		x"B3DA" when address_in = 16#0528# else
		x"C33D" when address_in = 16#0529# else
		x"D31C" when address_in = 16#052A# else
		x"E37F" when address_in = 16#052B# else
		x"F35E" when address_in = 16#052C# else
		x"02B1" when address_in = 16#052D# else
		x"1290" when address_in = 16#052E# else
		x"22F3" when address_in = 16#052F# else
		x"32D2" when address_in = 16#0530# else
		x"4235" when address_in = 16#0531# else
		x"5214" when address_in = 16#0532# else
		x"6277" when address_in = 16#0533# else
		x"7256" when address_in = 16#0534# else
		x"B5EA" when address_in = 16#0535# else
		x"A5CB" when address_in = 16#0536# else
		x"95A8" when address_in = 16#0537# else
		x"8589" when address_in = 16#0538# else
		x"F56E" when address_in = 16#0539# else
		x"E54F" when address_in = 16#053A# else
		x"D52C" when address_in = 16#053B# else
		x"C50D" when address_in = 16#053C# else
		x"34E2" when address_in = 16#053D# else
		x"24C3" when address_in = 16#053E# else
		x"14A0" when address_in = 16#053F# else
		x"0481" when address_in = 16#0540# else
		x"7466" when address_in = 16#0541# else
		x"6447" when address_in = 16#0542# else
		x"5424" when address_in = 16#0543# else
		x"4405" when address_in = 16#0544# else
		x"A7DB" when address_in = 16#0545# else
		x"B7FA" when address_in = 16#0546# else
		x"8799" when address_in = 16#0547# else
		x"97B8" when address_in = 16#0548# else
		x"E75F" when address_in = 16#0549# else
		x"F77E" when address_in = 16#054A# else
		x"C71D" when address_in = 16#054B# else
		x"D73C" when address_in = 16#054C# else
		x"26D3" when address_in = 16#054D# else
		x"36F2" when address_in = 16#054E# else
		x"0691" when address_in = 16#054F# else
		x"16B0" when address_in = 16#0550# else
		x"6657" when address_in = 16#0551# else
		x"7676" when address_in = 16#0552# else
		x"4615" when address_in = 16#0553# else
		x"5634" when address_in = 16#0554# else
		x"D94C" when address_in = 16#0555# else
		x"C96D" when address_in = 16#0556# else
		x"F90E" when address_in = 16#0557# else
		x"E92F" when address_in = 16#0558# else
		x"99C8" when address_in = 16#0559# else
		x"89E9" when address_in = 16#055A# else
		x"B98A" when address_in = 16#055B# else
		x"A9AB" when address_in = 16#055C# else
		x"5844" when address_in = 16#055D# else
		x"4865" when address_in = 16#055E# else
		x"7806" when address_in = 16#055F# else
		x"6827" when address_in = 16#0560# else
		x"18C0" when address_in = 16#0561# else
		x"08E1" when address_in = 16#0562# else
		x"3882" when address_in = 16#0563# else
		x"28A3" when address_in = 16#0564# else
		x"CB7D" when address_in = 16#0565# else
		x"DB5C" when address_in = 16#0566# else
		x"EB3F" when address_in = 16#0567# else
		x"FB1E" when address_in = 16#0568# else
		x"8BF9" when address_in = 16#0569# else
		x"9BD8" when address_in = 16#056A# else
		x"ABBB" when address_in = 16#056B# else
		x"BB9A" when address_in = 16#056C# else
		x"4A75" when address_in = 16#056D# else
		x"5A54" when address_in = 16#056E# else
		x"6A37" when address_in = 16#056F# else
		x"7A16" when address_in = 16#0570# else
		x"0AF1" when address_in = 16#0571# else
		x"1AD0" when address_in = 16#0572# else
		x"2AB3" when address_in = 16#0573# else
		x"3A92" when address_in = 16#0574# else
		x"FD2E" when address_in = 16#0575# else
		x"ED0F" when address_in = 16#0576# else
		x"DD6C" when address_in = 16#0577# else
		x"CD4D" when address_in = 16#0578# else
		x"BDAA" when address_in = 16#0579# else
		x"AD8B" when address_in = 16#057A# else
		x"9DE8" when address_in = 16#057B# else
		x"8DC9" when address_in = 16#057C# else
		x"7C26" when address_in = 16#057D# else
		x"6C07" when address_in = 16#057E# else
		x"5C64" when address_in = 16#057F# else
		x"4C45" when address_in = 16#0580# else
		x"3CA2" when address_in = 16#0581# else
		x"2C83" when address_in = 16#0582# else
		x"1CE0" when address_in = 16#0583# else
		x"0CC1" when address_in = 16#0584# else
		x"EF1F" when address_in = 16#0585# else
		x"FF3E" when address_in = 16#0586# else
		x"CF5D" when address_in = 16#0587# else
		x"DF7C" when address_in = 16#0588# else
		x"AF9B" when address_in = 16#0589# else
		x"BFBA" when address_in = 16#058A# else
		x"8FD9" when address_in = 16#058B# else
		x"9FF8" when address_in = 16#058C# else
		x"6E17" when address_in = 16#058D# else
		x"7E36" when address_in = 16#058E# else
		x"4E55" when address_in = 16#058F# else
		x"5E74" when address_in = 16#0590# else
		x"2E93" when address_in = 16#0591# else
		x"3EB2" when address_in = 16#0592# else
		x"0ED1" when address_in = 16#0593# else
		x"1EF0" when address_in = 16#0594# else
		x"2411" when address_in = 16#0595# else
		x"BE1F" when address_in = 16#0596# else
		x"EFCF" when address_in = 16#0597# else
		x"E0DF" when address_in = 16#0598# else
		x"BFDE" when address_in = 16#0599# else
		x"BFCD" when address_in = 16#059A# else
		x"E010" when address_in = 16#059B# else
		x"E6A0" when address_in = 16#059C# else
		x"E0B0" when address_in = 16#059D# else
		x"E4E8" when address_in = 16#059E# else
		x"E5FD" when address_in = 16#059F# else
		x"EF0F" when address_in = 16#05A0# else
		x"9503" when address_in = 16#05A1# else
		x"BF0B" when address_in = 16#05A2# else
		x"C004" when address_in = 16#05A3# else
		x"95D8" when address_in = 16#05A4# else
		x"920D" when address_in = 16#05A5# else
		x"9631" when address_in = 16#05A6# else
		x"F3C8" when address_in = 16#05A7# else
		x"37AA" when address_in = 16#05A8# else
		x"07B1" when address_in = 16#05A9# else
		x"F7C9" when address_in = 16#05AA# else
		x"E011" when address_in = 16#05AB# else
		x"E7AA" when address_in = 16#05AC# else
		x"E0B0" when address_in = 16#05AD# else
		x"C001" when address_in = 16#05AE# else
		x"921D" when address_in = 16#05AF# else
		x"37A6" when address_in = 16#05B0# else
		x"07B1" when address_in = 16#05B1# else
		x"F7E1" when address_in = 16#05B2# else
		x"940C" when address_in = 16#05B3# else
		x"05C6" when address_in = 16#05B4# else
		x"940C" when address_in = 16#05B5# else
		x"0000" when address_in = 16#05B6# else
		x"B38A" when address_in = 16#05B7# else
		x"6087" when address_in = 16#05B8# else
		x"BB8A" when address_in = 16#05B9# else
		x"9AD9" when address_in = 16#05BA# else
		x"9ADA" when address_in = 16#05BB# else
		x"9AD8" when address_in = 16#05BC# else
		x"E063" when address_in = 16#05BD# else
		x"E180" when address_in = 16#05BE# else
		x"940E" when address_in = 16#05BF# else
		x"2D62" when address_in = 16#05C0# else
		x"940E" when address_in = 16#05C1# else
		x"2C46" when address_in = 16#05C2# else
		x"940E" when address_in = 16#05C3# else
		x"25AF" when address_in = 16#05C4# else
		x"9508" when address_in = 16#05C5# else
		x"EFCF" when address_in = 16#05C6# else
		x"E0DF" when address_in = 16#05C7# else
		x"BFDE" when address_in = 16#05C8# else
		x"BFCD" when address_in = 16#05C9# else
		x"E080" when address_in = 16#05CA# else
		x"940E" when address_in = 16#05CB# else
		x"05D1" when address_in = 16#05CC# else
		x"E080" when address_in = 16#05CD# else
		x"E090" when address_in = 16#05CE# else
		x"940C" when address_in = 16#05CF# else
		x"2EA3" when address_in = 16#05D0# else
		x"931F" when address_in = 16#05D1# else
		x"2F18" when address_in = 16#05D2# else
		x"94F8" when address_in = 16#05D3# else
		x"940E" when address_in = 16#05D4# else
		x"2D93" when address_in = 16#05D5# else
		x"940E" when address_in = 16#05D6# else
		x"242B" when address_in = 16#05D7# else
		x"940E" when address_in = 16#05D8# else
		x"0979" when address_in = 16#05D9# else
		x"940E" when address_in = 16#05DA# else
		x"1164" when address_in = 16#05DB# else
		x"940E" when address_in = 16#05DC# else
		x"2568" when address_in = 16#05DD# else
		x"2F81" when address_in = 16#05DE# else
		x"940E" when address_in = 16#05DF# else
		x"0BF3" when address_in = 16#05E0# else
		x"940E" when address_in = 16#05E1# else
		x"1541" when address_in = 16#05E2# else
		x"940E" when address_in = 16#05E3# else
		x"22B5" when address_in = 16#05E4# else
		x"940E" when address_in = 16#05E5# else
		x"05B7" when address_in = 16#05E6# else
		x"9478" when address_in = 16#05E7# else
		x"940E" when address_in = 16#05E8# else
		x"0B0A" when address_in = 16#05E9# else
		x"940E" when address_in = 16#05EA# else
		x"0F1A" when address_in = 16#05EB# else
		x"E080" when address_in = 16#05EC# else
		x"E090" when address_in = 16#05ED# else
		x"911F" when address_in = 16#05EE# else
		x"9508" when address_in = 16#05EF# else
		x"2FB9" when address_in = 16#05F0# else
		x"2FA8" when address_in = 16#05F1# else
		x"2FF7" when address_in = 16#05F2# else
		x"2FE6" when address_in = 16#05F3# else
		x"8186" when address_in = 16#05F4# else
		x"2799" when address_in = 16#05F5# else
		x"3082" when address_in = 16#05F6# else
		x"0591" when address_in = 16#05F7# else
		x"F0F1" when address_in = 16#05F8# else
		x"3083" when address_in = 16#05F9# else
		x"0591" when address_in = 16#05FA# else
		x"F41C" when address_in = 16#05FB# else
		x"2B89" when address_in = 16#05FC# else
		x"F021" when address_in = 16#05FD# else
		x"C01C" when address_in = 16#05FE# else
		x"9706" when address_in = 16#05FF# else
		x"F091" when address_in = 16#0600# else
		x"C019" when address_in = 16#0601# else
		x"8180" when address_in = 16#0602# else
		x"938C" when address_in = 16#0603# else
		x"2FFB" when address_in = 16#0604# else
		x"2FEA" when address_in = 16#0605# else
		x"8211" when address_in = 16#0606# else
		x"E087" when address_in = 16#0607# else
		x"940E" when address_in = 16#0608# else
		x"0420" when address_in = 16#0609# else
		x"E020" when address_in = 16#060A# else
		x"E144" when address_in = 16#060B# else
		x"E050" when address_in = 16#060C# else
		x"E060" when address_in = 16#060D# else
		x"E070" when address_in = 16#060E# else
		x"2F82" when address_in = 16#060F# else
		x"940E" when address_in = 16#0610# else
		x"040A" when address_in = 16#0611# else
		x"C00B" when address_in = 16#0612# else
		x"E080" when address_in = 16#0613# else
		x"940E" when address_in = 16#0614# else
		x"040E" when address_in = 16#0615# else
		x"C007" when address_in = 16#0616# else
		x"E088" when address_in = 16#0617# else
		x"940E" when address_in = 16#0618# else
		x"0420" when address_in = 16#0619# else
		x"C003" when address_in = 16#061A# else
		x"EE8A" when address_in = 16#061B# else
		x"EF9F" when address_in = 16#061C# else
		x"9508" when address_in = 16#061D# else
		x"E080" when address_in = 16#061E# else
		x"E090" when address_in = 16#061F# else
		x"9508" when address_in = 16#0620# else
		x"E080" when address_in = 16#0621# else
		x"E099" when address_in = 16#0622# else
		x"27AA" when address_in = 16#0623# else
		x"FD97" when address_in = 16#0624# else
		x"95A0" when address_in = 16#0625# else
		x"2FBA" when address_in = 16#0626# else
		x"95B6" when address_in = 16#0627# else
		x"95A7" when address_in = 16#0628# else
		x"9597" when address_in = 16#0629# else
		x"9587" when address_in = 16#062A# else
		x"9508" when address_in = 16#062B# else
		x"93CF" when address_in = 16#062C# else
		x"93DF" when address_in = 16#062D# else
		x"2FF9" when address_in = 16#062E# else
		x"2FE8" when address_in = 16#062F# else
		x"81A3" when address_in = 16#0630# else
		x"81B4" when address_in = 16#0631# else
		x"8185" when address_in = 16#0632# else
		x"8196" when address_in = 16#0633# else
		x"2FDB" when address_in = 16#0634# else
		x"2FCA" when address_in = 16#0635# else
		x"839E" when address_in = 16#0636# else
		x"838D" when address_in = 16#0637# else
		x"8005" when address_in = 16#0638# else
		x"81F6" when address_in = 16#0639# else
		x"2DE0" when address_in = 16#063A# else
		x"83B4" when address_in = 16#063B# else
		x"83A3" when address_in = 16#063C# else
		x"91DF" when address_in = 16#063D# else
		x"91CF" when address_in = 16#063E# else
		x"9508" when address_in = 16#063F# else
		x"92AF" when address_in = 16#0640# else
		x"92BF" when address_in = 16#0641# else
		x"92CF" when address_in = 16#0642# else
		x"92DF" when address_in = 16#0643# else
		x"92EF" when address_in = 16#0644# else
		x"92FF" when address_in = 16#0645# else
		x"930F" when address_in = 16#0646# else
		x"931F" when address_in = 16#0647# else
		x"93CF" when address_in = 16#0648# else
		x"93DF" when address_in = 16#0649# else
		x"2EA6" when address_in = 16#064A# else
		x"24CC" when address_in = 16#064B# else
		x"24DD" when address_in = 16#064C# else
		x"9700" when address_in = 16#064D# else
		x"F419" when address_in = 16#064E# else
		x"2D9D" when address_in = 16#064F# else
		x"2D8C" when address_in = 16#0650# else
		x"C0A3" when address_in = 16#0651# else
		x"E05A" when address_in = 16#0652# else
		x"2EE5" when address_in = 16#0653# else
		x"2CF1" when address_in = 16#0654# else
		x"0EE8" when address_in = 16#0655# else
		x"1EF9" when address_in = 16#0656# else
		x"E043" when address_in = 16#0657# else
		x"94F6" when address_in = 16#0658# else
		x"94E7" when address_in = 16#0659# else
		x"954A" when address_in = 16#065A# else
		x"F7E1" when address_in = 16#065B# else
		x"B6BF" when address_in = 16#065C# else
		x"94F8" when address_in = 16#065D# else
		x"91E0" when address_in = 16#065E# else
		x"007C" when address_in = 16#065F# else
		x"91F0" when address_in = 16#0660# else
		x"007D" when address_in = 16#0661# else
		x"81C5" when address_in = 16#0662# else
		x"81D6" when address_in = 16#0663# else
		x"17CE" when address_in = 16#0664# else
		x"07DF" when address_in = 16#0665# else
		x"F141" when address_in = 16#0666# else
		x"8108" when address_in = 16#0667# else
		x"8119" when address_in = 16#0668# else
		x"E033" when address_in = 16#0669# else
		x"0F00" when address_in = 16#066A# else
		x"1F11" when address_in = 16#066B# else
		x"953A" when address_in = 16#066C# else
		x"F7E1" when address_in = 16#066D# else
		x"0F0C" when address_in = 16#066E# else
		x"1F1D" when address_in = 16#066F# else
		x"2FF1" when address_in = 16#0670# else
		x"2FE0" when address_in = 16#0671# else
		x"8180" when address_in = 16#0672# else
		x"8191" when address_in = 16#0673# else
		x"2399" when address_in = 16#0674# else
		x"F07C" when address_in = 16#0675# else
		x"2F91" when address_in = 16#0676# else
		x"2F80" when address_in = 16#0677# else
		x"940E" when address_in = 16#0678# else
		x"062C" when address_in = 16#0679# else
		x"8188" when address_in = 16#067A# else
		x"8199" when address_in = 16#067B# else
		x"2FF1" when address_in = 16#067C# else
		x"2FE0" when address_in = 16#067D# else
		x"8120" when address_in = 16#067E# else
		x"8131" when address_in = 16#067F# else
		x"0F82" when address_in = 16#0680# else
		x"1F93" when address_in = 16#0681# else
		x"8399" when address_in = 16#0682# else
		x"8388" when address_in = 16#0683# else
		x"CFE2" when address_in = 16#0684# else
		x"800D" when address_in = 16#0685# else
		x"81DE" when address_in = 16#0686# else
		x"2DC0" when address_in = 16#0687# else
		x"9180" when address_in = 16#0688# else
		x"007C" when address_in = 16#0689# else
		x"9190" when address_in = 16#068A# else
		x"007D" when address_in = 16#068B# else
		x"17C8" when address_in = 16#068C# else
		x"07D9" when address_in = 16#068D# else
		x"F6C1" when address_in = 16#068E# else
		x"91E0" when address_in = 16#068F# else
		x"007C" when address_in = 16#0690# else
		x"91F0" when address_in = 16#0691# else
		x"007D" when address_in = 16#0692# else
		x"81C5" when address_in = 16#0693# else
		x"81D6" when address_in = 16#0694# else
		x"17CE" when address_in = 16#0695# else
		x"07DF" when address_in = 16#0696# else
		x"F099" when address_in = 16#0697# else
		x"16CC" when address_in = 16#0698# else
		x"06DD" when address_in = 16#0699# else
		x"F438" when address_in = 16#069A# else
		x"8188" when address_in = 16#069B# else
		x"8199" when address_in = 16#069C# else
		x"158E" when address_in = 16#069D# else
		x"059F" when address_in = 16#069E# else
		x"F010" when address_in = 16#069F# else
		x"2ECC" when address_in = 16#06A0# else
		x"2EDD" when address_in = 16#06A1# else
		x"800D" when address_in = 16#06A2# else
		x"81DE" when address_in = 16#06A3# else
		x"2DC0" when address_in = 16#06A4# else
		x"17CE" when address_in = 16#06A5# else
		x"07DF" when address_in = 16#06A6# else
		x"F781" when address_in = 16#06A7# else
		x"14C1" when address_in = 16#06A8# else
		x"04D1" when address_in = 16#06A9# else
		x"F421" when address_in = 16#06AA# else
		x"BEBF" when address_in = 16#06AB# else
		x"E080" when address_in = 16#06AC# else
		x"E090" when address_in = 16#06AD# else
		x"C046" when address_in = 16#06AE# else
		x"2DFD" when address_in = 16#06AF# else
		x"2DEC" when address_in = 16#06B0# else
		x"8180" when address_in = 16#06B1# else
		x"8191" when address_in = 16#06B2# else
		x"198E" when address_in = 16#06B3# else
		x"099F" when address_in = 16#06B4# else
		x"2FD9" when address_in = 16#06B5# else
		x"2FC8" when address_in = 16#06B6# else
		x"E023" when address_in = 16#06B7# else
		x"0FCC" when address_in = 16#06B8# else
		x"1FDD" when address_in = 16#06B9# else
		x"952A" when address_in = 16#06BA# else
		x"F7E1" when address_in = 16#06BB# else
		x"0DCC" when address_in = 16#06BC# else
		x"1DDD" when address_in = 16#06BD# else
		x"15CC" when address_in = 16#06BE# else
		x"05DD" when address_in = 16#06BF# else
		x"F429" when address_in = 16#06C0# else
		x"2F8C" when address_in = 16#06C1# else
		x"2F9D" when address_in = 16#06C2# else
		x"940E" when address_in = 16#06C3# else
		x"062C" when address_in = 16#06C4# else
		x"C006" when address_in = 16#06C5# else
		x"2DFD" when address_in = 16#06C6# else
		x"2DEC" when address_in = 16#06C7# else
		x"8391" when address_in = 16#06C8# else
		x"8380" when address_in = 16#06C9# else
		x"82F9" when address_in = 16#06CA# else
		x"82E8" when address_in = 16#06CB# else
		x"8188" when address_in = 16#06CC# else
		x"8199" when address_in = 16#06CD# else
		x"6890" when address_in = 16#06CE# else
		x"8399" when address_in = 16#06CF# else
		x"8388" when address_in = 16#06D0# else
		x"82AA" when address_in = 16#06D1# else
		x"2D8A" when address_in = 16#06D2# else
		x"940E" when address_in = 16#06D3# else
		x"2D9E" when address_in = 16#06D4# else
		x"2F18" when address_in = 16#06D5# else
		x"7017" when address_in = 16#06D6# else
		x"2F81" when address_in = 16#06D7# else
		x"6088" when address_in = 16#06D8# else
		x"2F48" when address_in = 16#06D9# else
		x"E068" when address_in = 16#06DA# else
		x"E070" when address_in = 16#06DB# else
		x"2F8C" when address_in = 16#06DC# else
		x"2F9D" when address_in = 16#06DD# else
		x"940E" when address_in = 16#06DE# else
		x"0A4B" when address_in = 16#06DF# else
		x"E083" when address_in = 16#06E0# else
		x"0CEE" when address_in = 16#06E1# else
		x"1CFF" when address_in = 16#06E2# else
		x"958A" when address_in = 16#06E3# else
		x"F7E1" when address_in = 16#06E4# else
		x"EF88" when address_in = 16#06E5# else
		x"EF9F" when address_in = 16#06E6# else
		x"0EE8" when address_in = 16#06E7# else
		x"1EF9" when address_in = 16#06E8# else
		x"2F41" when address_in = 16#06E9# else
		x"2D7F" when address_in = 16#06EA# else
		x"2D6E" when address_in = 16#06EB# else
		x"2F8C" when address_in = 16#06EC# else
		x"2F9D" when address_in = 16#06ED# else
		x"9608" when address_in = 16#06EE# else
		x"940E" when address_in = 16#06EF# else
		x"0A4B" when address_in = 16#06F0# else
		x"BEBF" when address_in = 16#06F1# else
		x"2F8C" when address_in = 16#06F2# else
		x"2F9D" when address_in = 16#06F3# else
		x"9603" when address_in = 16#06F4# else
		x"91DF" when address_in = 16#06F5# else
		x"91CF" when address_in = 16#06F6# else
		x"911F" when address_in = 16#06F7# else
		x"910F" when address_in = 16#06F8# else
		x"90FF" when address_in = 16#06F9# else
		x"90EF" when address_in = 16#06FA# else
		x"90DF" when address_in = 16#06FB# else
		x"90CF" when address_in = 16#06FC# else
		x"90BF" when address_in = 16#06FD# else
		x"90AF" when address_in = 16#06FE# else
		x"9508" when address_in = 16#06FF# else
		x"925F" when address_in = 16#0700# else
		x"926F" when address_in = 16#0701# else
		x"927F" when address_in = 16#0702# else
		x"928F" when address_in = 16#0703# else
		x"929F" when address_in = 16#0704# else
		x"92AF" when address_in = 16#0705# else
		x"92BF" when address_in = 16#0706# else
		x"92CF" when address_in = 16#0707# else
		x"92DF" when address_in = 16#0708# else
		x"92EF" when address_in = 16#0709# else
		x"92FF" when address_in = 16#070A# else
		x"930F" when address_in = 16#070B# else
		x"931F" when address_in = 16#070C# else
		x"93CF" when address_in = 16#070D# else
		x"93DF" when address_in = 16#070E# else
		x"B7CD" when address_in = 16#070F# else
		x"B7DE" when address_in = 16#0710# else
		x"9726" when address_in = 16#0711# else
		x"B60F" when address_in = 16#0712# else
		x"94F8" when address_in = 16#0713# else
		x"BFDE" when address_in = 16#0714# else
		x"BE0F" when address_in = 16#0715# else
		x"BFCD" when address_in = 16#0716# else
		x"2E68" when address_in = 16#0717# else
		x"2E79" when address_in = 16#0718# else
		x"2E56" when address_in = 16#0719# else
		x"8349" when address_in = 16#071A# else
		x"9703" when address_in = 16#071B# else
		x"839B" when address_in = 16#071C# else
		x"838A" when address_in = 16#071D# else
		x"EF9F" when address_in = 16#071E# else
		x"1769" when address_in = 16#071F# else
		x"F409" when address_in = 16#0720# else
		x"C092" when address_in = 16#0721# else
		x"1461" when address_in = 16#0722# else
		x"0471" when address_in = 16#0723# else
		x"F409" when address_in = 16#0724# else
		x"C08E" when address_in = 16#0725# else
		x"B6EF" when address_in = 16#0726# else
		x"94F8" when address_in = 16#0727# else
		x"9180" when address_in = 16#0728# else
		x"0171" when address_in = 16#0729# else
		x"9190" when address_in = 16#072A# else
		x"0172" when address_in = 16#072B# else
		x"80CA" when address_in = 16#072C# else
		x"80DB" when address_in = 16#072D# else
		x"1AC8" when address_in = 16#072E# else
		x"0AD9" when address_in = 16#072F# else
		x"2DFD" when address_in = 16#0730# else
		x"2DEC" when address_in = 16#0731# else
		x"E0A4" when address_in = 16#0732# else
		x"95F6" when address_in = 16#0733# else
		x"95E7" when address_in = 16#0734# else
		x"95AA" when address_in = 16#0735# else
		x"F7E1" when address_in = 16#0736# else
		x"83FD" when address_in = 16#0737# else
		x"83EC" when address_in = 16#0738# else
		x"2D1D" when address_in = 16#0739# else
		x"2D0C" when address_in = 16#073A# else
		x"9516" when address_in = 16#073B# else
		x"9507" when address_in = 16#073C# else
		x"2E8E" when address_in = 16#073D# else
		x"2E9F" when address_in = 16#073E# else
		x"E980" when address_in = 16#073F# else
		x"E099" when address_in = 16#0740# else
		x"0E88" when address_in = 16#0741# else
		x"1E99" when address_in = 16#0742# else
		x"2DF9" when address_in = 16#0743# else
		x"2DE8" when address_in = 16#0744# else
		x"80F0" when address_in = 16#0745# else
		x"2D8F" when address_in = 16#0746# else
		x"2799" when address_in = 16#0747# else
		x"7004" when address_in = 16#0748# else
		x"7010" when address_in = 16#0749# else
		x"2E00" when address_in = 16#074A# else
		x"C002" when address_in = 16#074B# else
		x"9595" when address_in = 16#074C# else
		x"9587" when address_in = 16#074D# else
		x"940A" when address_in = 16#074E# else
		x"F7E2" when address_in = 16#074F# else
		x"2EF8" when address_in = 16#0750# else
		x"E0FF" when address_in = 16#0751# else
		x"22FF" when address_in = 16#0752# else
		x"2CAF" when address_in = 16#0753# else
		x"24BB" when address_in = 16#0754# else
		x"2D9B" when address_in = 16#0755# else
		x"2D8A" when address_in = 16#0756# else
		x"7088" when address_in = 16#0757# else
		x"7090" when address_in = 16#0758# else
		x"5F87" when address_in = 16#0759# else
		x"4F9F" when address_in = 16#075A# else
		x"F421" when address_in = 16#075B# else
		x"BEEF" when address_in = 16#075C# else
		x"E085" when address_in = 16#075D# else
		x"940E" when address_in = 16#075E# else
		x"2E07" when address_in = 16#075F# else
		x"E087" when address_in = 16#0760# else
		x"22A8" when address_in = 16#0761# else
		x"24BB" when address_in = 16#0762# else
		x"81E9" when address_in = 16#0763# else
		x"2F8E" when address_in = 16#0764# else
		x"2799" when address_in = 16#0765# else
		x"16A8" when address_in = 16#0766# else
		x"06B9" when address_in = 16#0767# else
		x"F019" when address_in = 16#0768# else
		x"30E7" when address_in = 16#0769# else
		x"F009" when address_in = 16#076A# else
		x"C044" when address_in = 16#076B# else
		x"2D85" when address_in = 16#076C# else
		x"940E" when address_in = 16#076D# else
		x"2D9E" when address_in = 16#076E# else
		x"838E" when address_in = 16#076F# else
		x"FF87" when address_in = 16#0770# else
		x"C004" when address_in = 16#0771# else
		x"BEEF" when address_in = 16#0772# else
		x"E086" when address_in = 16#0773# else
		x"940E" when address_in = 16#0774# else
		x"2E07" when address_in = 16#0775# else
		x"81FE" when address_in = 16#0776# else
		x"2F4F" when address_in = 16#0777# else
		x"2755" when address_in = 16#0778# else
		x"FD47" when address_in = 16#0779# else
		x"9550" when address_in = 16#077A# else
		x"154A" when address_in = 16#077B# else
		x"055B" when address_in = 16#077C# else
		x"F1C9" when address_in = 16#077D# else
		x"2DF9" when address_in = 16#077E# else
		x"2DE8" when address_in = 16#077F# else
		x"8120" when address_in = 16#0780# else
		x"E08F" when address_in = 16#0781# else
		x"E090" when address_in = 16#0782# else
		x"2E00" when address_in = 16#0783# else
		x"C002" when address_in = 16#0784# else
		x"0F88" when address_in = 16#0785# else
		x"1F99" when address_in = 16#0786# else
		x"940A" when address_in = 16#0787# else
		x"F7E2" when address_in = 16#0788# else
		x"9580" when address_in = 16#0789# else
		x"2328" when address_in = 16#078A# else
		x"7047" when address_in = 16#078B# else
		x"7050" when address_in = 16#078C# else
		x"6048" when address_in = 16#078D# else
		x"C002" when address_in = 16#078E# else
		x"0F44" when address_in = 16#078F# else
		x"1F55" when address_in = 16#0790# else
		x"950A" when address_in = 16#0791# else
		x"F7E2" when address_in = 16#0792# else
		x"2B24" when address_in = 16#0793# else
		x"EC8C" when address_in = 16#0794# else
		x"BB8B" when address_in = 16#0795# else
		x"BB2B" when address_in = 16#0796# else
		x"81FC" when address_in = 16#0797# else
		x"BBFB" when address_in = 16#0798# else
		x"2CCD" when address_in = 16#0799# else
		x"24DD" when address_in = 16#079A# else
		x"94C2" when address_in = 16#079B# else
		x"E06F" when address_in = 16#079C# else
		x"22C6" when address_in = 16#079D# else
		x"BACB" when address_in = 16#079E# else
		x"2DF9" when address_in = 16#079F# else
		x"2DE8" when address_in = 16#07A0# else
		x"8320" when address_in = 16#07A1# else
		x"81FE" when address_in = 16#07A2# else
		x"70F7" when address_in = 16#07A3# else
		x"83FE" when address_in = 16#07A4# else
		x"E027" when address_in = 16#07A5# else
		x"22F2" when address_in = 16#07A6# else
		x"2F2F" when address_in = 16#07A7# else
		x"2D4F" when address_in = 16#07A8# else
		x"E06F" when address_in = 16#07A9# else
		x"2D97" when address_in = 16#07AA# else
		x"2D86" when address_in = 16#07AB# else
		x"9605" when address_in = 16#07AC# else
		x"940E" when address_in = 16#07AD# else
		x"0AA0" when address_in = 16#07AE# else
		x"C007" when address_in = 16#07AF# else
		x"BEEF" when address_in = 16#07B0# else
		x"E085" when address_in = 16#07B1# else
		x"940E" when address_in = 16#07B2# else
		x"2E07" when address_in = 16#07B3# else
		x"EE8A" when address_in = 16#07B4# else
		x"EF9F" when address_in = 16#07B5# else
		x"C006" when address_in = 16#07B6# else
		x"BEEF" when address_in = 16#07B7# else
		x"81EA" when address_in = 16#07B8# else
		x"81FB" when address_in = 16#07B9# else
		x"8252" when address_in = 16#07BA# else
		x"E080" when address_in = 16#07BB# else
		x"E090" when address_in = 16#07BC# else
		x"9626" when address_in = 16#07BD# else
		x"B60F" when address_in = 16#07BE# else
		x"94F8" when address_in = 16#07BF# else
		x"BFDE" when address_in = 16#07C0# else
		x"BE0F" when address_in = 16#07C1# else
		x"BFCD" when address_in = 16#07C2# else
		x"91DF" when address_in = 16#07C3# else
		x"91CF" when address_in = 16#07C4# else
		x"911F" when address_in = 16#07C5# else
		x"910F" when address_in = 16#07C6# else
		x"90FF" when address_in = 16#07C7# else
		x"90EF" when address_in = 16#07C8# else
		x"90DF" when address_in = 16#07C9# else
		x"90CF" when address_in = 16#07CA# else
		x"90BF" when address_in = 16#07CB# else
		x"90AF" when address_in = 16#07CC# else
		x"909F" when address_in = 16#07CD# else
		x"908F" when address_in = 16#07CE# else
		x"907F" when address_in = 16#07CF# else
		x"906F" when address_in = 16#07D0# else
		x"905F" when address_in = 16#07D1# else
		x"9508" when address_in = 16#07D2# else
		x"93CF" when address_in = 16#07D3# else
		x"93DF" when address_in = 16#07D4# else
		x"2FF9" when address_in = 16#07D5# else
		x"2FE8" when address_in = 16#07D6# else
		x"91A0" when address_in = 16#07D7# else
		x"007C" when address_in = 16#07D8# else
		x"91B0" when address_in = 16#07D9# else
		x"007D" when address_in = 16#07DA# else
		x"2FDB" when address_in = 16#07DB# else
		x"2FCA" when address_in = 16#07DC# else
		x"818D" when address_in = 16#07DD# else
		x"819E" when address_in = 16#07DE# else
		x"83FE" when address_in = 16#07DF# else
		x"83ED" when address_in = 16#07E0# else
		x"83B4" when address_in = 16#07E1# else
		x"83A3" when address_in = 16#07E2# else
		x"8396" when address_in = 16#07E3# else
		x"8385" when address_in = 16#07E4# else
		x"2FD9" when address_in = 16#07E5# else
		x"2FC8" when address_in = 16#07E6# else
		x"83FC" when address_in = 16#07E7# else
		x"83EB" when address_in = 16#07E8# else
		x"91DF" when address_in = 16#07E9# else
		x"91CF" when address_in = 16#07EA# else
		x"9508" when address_in = 16#07EB# else
		x"931F" when address_in = 16#07EC# else
		x"93CF" when address_in = 16#07ED# else
		x"93DF" when address_in = 16#07EE# else
		x"9700" when address_in = 16#07EF# else
		x"F409" when address_in = 16#07F0# else
		x"C093" when address_in = 16#07F1# else
		x"2FD9" when address_in = 16#07F2# else
		x"2FC8" when address_in = 16#07F3# else
		x"9723" when address_in = 16#07F4# else
		x"E041" when address_in = 16#07F5# else
		x"39C0" when address_in = 16#07F6# else
		x"07D4" when address_in = 16#07F7# else
		x"F408" when address_in = 16#07F8# else
		x"C08B" when address_in = 16#07F9# else
		x"9180" when address_in = 16#07FA# else
		x"007E" when address_in = 16#07FB# else
		x"9190" when address_in = 16#07FC# else
		x"007F" when address_in = 16#07FD# else
		x"E0E3" when address_in = 16#07FE# else
		x"0F88" when address_in = 16#07FF# else
		x"1F99" when address_in = 16#0800# else
		x"95EA" when address_in = 16#0801# else
		x"F7E1" when address_in = 16#0802# else
		x"5780" when address_in = 16#0803# else
		x"4F9E" when address_in = 16#0804# else
		x"17C8" when address_in = 16#0805# else
		x"07D9" when address_in = 16#0806# else
		x"F008" when address_in = 16#0807# else
		x"C07C" when address_in = 16#0808# else
		x"B71F" when address_in = 16#0809# else
		x"94F8" when address_in = 16#080A# else
		x"9180" when address_in = 16#080B# else
		x"0171" when address_in = 16#080C# else
		x"9190" when address_in = 16#080D# else
		x"0172" when address_in = 16#080E# else
		x"2FFD" when address_in = 16#080F# else
		x"2FEC" when address_in = 16#0810# else
		x"1BE8" when address_in = 16#0811# else
		x"0BF9" when address_in = 16#0812# else
		x"2FAE" when address_in = 16#0813# else
		x"2FBF" when address_in = 16#0814# else
		x"E073" when address_in = 16#0815# else
		x"95B6" when address_in = 16#0816# else
		x"95A7" when address_in = 16#0817# else
		x"957A" when address_in = 16#0818# else
		x"F7E1" when address_in = 16#0819# else
		x"E054" when address_in = 16#081A# else
		x"95F6" when address_in = 16#081B# else
		x"95E7" when address_in = 16#081C# else
		x"955A" when address_in = 16#081D# else
		x"F7E1" when address_in = 16#081E# else
		x"2F2A" when address_in = 16#081F# else
		x"2F3B" when address_in = 16#0820# else
		x"7021" when address_in = 16#0821# else
		x"7030" when address_in = 16#0822# else
		x"57E0" when address_in = 16#0823# else
		x"4FF6" when address_in = 16#0824# else
		x"8150" when address_in = 16#0825# else
		x"2F85" when address_in = 16#0826# else
		x"2799" when address_in = 16#0827# else
		x"0F22" when address_in = 16#0828# else
		x"1F33" when address_in = 16#0829# else
		x"0F22" when address_in = 16#082A# else
		x"1F33" when address_in = 16#082B# else
		x"C002" when address_in = 16#082C# else
		x"9595" when address_in = 16#082D# else
		x"9587" when address_in = 16#082E# else
		x"952A" when address_in = 16#082F# else
		x"F7E2" when address_in = 16#0830# else
		x"2F58" when address_in = 16#0831# else
		x"705F" when address_in = 16#0832# else
		x"2F25" when address_in = 16#0833# else
		x"2733" when address_in = 16#0834# else
		x"2F93" when address_in = 16#0835# else
		x"2F82" when address_in = 16#0836# else
		x"7088" when address_in = 16#0837# else
		x"7090" when address_in = 16#0838# else
		x"5F87" when address_in = 16#0839# else
		x"4F9F" when address_in = 16#083A# else
		x"F411" when address_in = 16#083B# else
		x"BF1F" when address_in = 16#083C# else
		x"C00A" when address_in = 16#083D# else
		x"3067" when address_in = 16#083E# else
		x"F061" when address_in = 16#083F# else
		x"7027" when address_in = 16#0840# else
		x"7030" when address_in = 16#0841# else
		x"2F86" when address_in = 16#0842# else
		x"2799" when address_in = 16#0843# else
		x"1728" when address_in = 16#0844# else
		x"0739" when address_in = 16#0845# else
		x"F029" when address_in = 16#0846# else
		x"BF1F" when address_in = 16#0847# else
		x"E085" when address_in = 16#0848# else
		x"940E" when address_in = 16#0849# else
		x"2E07" when address_in = 16#084A# else
		x"C039" when address_in = 16#084B# else
		x"B71F" when address_in = 16#084C# else
		x"94F8" when address_in = 16#084D# else
		x"8188" when address_in = 16#084E# else
		x"8199" when address_in = 16#084F# else
		x"779F" when address_in = 16#0850# else
		x"8399" when address_in = 16#0851# else
		x"8388" when address_in = 16#0852# else
		x"EF8F" when address_in = 16#0853# else
		x"838A" when address_in = 16#0854# else
		x"2F6A" when address_in = 16#0855# else
		x"2F7B" when address_in = 16#0856# else
		x"9576" when address_in = 16#0857# else
		x"9567" when address_in = 16#0858# else
		x"2F2A" when address_in = 16#0859# else
		x"2F3B" when address_in = 16#085A# else
		x"7021" when address_in = 16#085B# else
		x"7030" when address_in = 16#085C# else
		x"2FF7" when address_in = 16#085D# else
		x"2FE6" when address_in = 16#085E# else
		x"57E0" when address_in = 16#085F# else
		x"4FF6" when address_in = 16#0860# else
		x"8140" when address_in = 16#0861# else
		x"0F22" when address_in = 16#0862# else
		x"1F33" when address_in = 16#0863# else
		x"0F22" when address_in = 16#0864# else
		x"1F33" when address_in = 16#0865# else
		x"E08F" when address_in = 16#0866# else
		x"E090" when address_in = 16#0867# else
		x"C002" when address_in = 16#0868# else
		x"0F88" when address_in = 16#0869# else
		x"1F99" when address_in = 16#086A# else
		x"952A" when address_in = 16#086B# else
		x"F7E2" when address_in = 16#086C# else
		x"2B48" when address_in = 16#086D# else
		x"EC8C" when address_in = 16#086E# else
		x"BB8B" when address_in = 16#086F# else
		x"BB4B" when address_in = 16#0870# else
		x"BB6B" when address_in = 16#0871# else
		x"2FAB" when address_in = 16#0872# else
		x"27BB" when address_in = 16#0873# else
		x"95A6" when address_in = 16#0874# else
		x"BBAB" when address_in = 16#0875# else
		x"8340" when address_in = 16#0876# else
		x"7057" when address_in = 16#0877# else
		x"E02F" when address_in = 16#0878# else
		x"2F45" when address_in = 16#0879# else
		x"2F62" when address_in = 16#087A# else
		x"2F8C" when address_in = 16#087B# else
		x"2F9D" when address_in = 16#087C# else
		x"9608" when address_in = 16#087D# else
		x"940E" when address_in = 16#087E# else
		x"0AA0" when address_in = 16#087F# else
		x"2F8C" when address_in = 16#0880# else
		x"2F9D" when address_in = 16#0881# else
		x"940E" when address_in = 16#0882# else
		x"07D3" when address_in = 16#0883# else
		x"BF1F" when address_in = 16#0884# else
		x"91DF" when address_in = 16#0885# else
		x"91CF" when address_in = 16#0886# else
		x"911F" when address_in = 16#0887# else
		x"9508" when address_in = 16#0888# else
		x"92BF" when address_in = 16#0889# else
		x"92CF" when address_in = 16#088A# else
		x"92DF" when address_in = 16#088B# else
		x"92EF" when address_in = 16#088C# else
		x"92FF" when address_in = 16#088D# else
		x"930F" when address_in = 16#088E# else
		x"931F" when address_in = 16#088F# else
		x"93CF" when address_in = 16#0890# else
		x"93DF" when address_in = 16#0891# else
		x"2EB6" when address_in = 16#0892# else
		x"2F14" when address_in = 16#0893# else
		x"9700" when address_in = 16#0894# else
		x"F409" when address_in = 16#0895# else
		x"C0A1" when address_in = 16#0896# else
		x"E02A" when address_in = 16#0897# else
		x"2EC2" when address_in = 16#0898# else
		x"2CD1" when address_in = 16#0899# else
		x"0EC8" when address_in = 16#089A# else
		x"1ED9" when address_in = 16#089B# else
		x"E093" when address_in = 16#089C# else
		x"94D6" when address_in = 16#089D# else
		x"94C7" when address_in = 16#089E# else
		x"959A" when address_in = 16#089F# else
		x"F7E1" when address_in = 16#08A0# else
		x"B70F" when address_in = 16#08A1# else
		x"94F8" when address_in = 16#08A2# else
		x"91E0" when address_in = 16#08A3# else
		x"007C" when address_in = 16#08A4# else
		x"91F0" when address_in = 16#08A5# else
		x"007D" when address_in = 16#08A6# else
		x"80E5" when address_in = 16#08A7# else
		x"80F6" when address_in = 16#08A8# else
		x"16EE" when address_in = 16#08A9# else
		x"06FF" when address_in = 16#08AA# else
		x"F191" when address_in = 16#08AB# else
		x"2DBF" when address_in = 16#08AC# else
		x"2DAE" when address_in = 16#08AD# else
		x"91CD" when address_in = 16#08AE# else
		x"91DC" when address_in = 16#08AF# else
		x"E083" when address_in = 16#08B0# else
		x"0FCC" when address_in = 16#08B1# else
		x"1FDD" when address_in = 16#08B2# else
		x"958A" when address_in = 16#08B3# else
		x"F7E1" when address_in = 16#08B4# else
		x"0DCE" when address_in = 16#08B5# else
		x"1DDF" when address_in = 16#08B6# else
		x"8188" when address_in = 16#08B7# else
		x"8199" when address_in = 16#08B8# else
		x"2399" when address_in = 16#08B9# else
		x"F08C" when address_in = 16#08BA# else
		x"2F8C" when address_in = 16#08BB# else
		x"2F9D" when address_in = 16#08BC# else
		x"940E" when address_in = 16#08BD# else
		x"062C" when address_in = 16#08BE# else
		x"2DFF" when address_in = 16#08BF# else
		x"2DEE" when address_in = 16#08C0# else
		x"8180" when address_in = 16#08C1# else
		x"8191" when address_in = 16#08C2# else
		x"8128" when address_in = 16#08C3# else
		x"8139" when address_in = 16#08C4# else
		x"0F82" when address_in = 16#08C5# else
		x"1F93" when address_in = 16#08C6# else
		x"8391" when address_in = 16#08C7# else
		x"8380" when address_in = 16#08C8# else
		x"158C" when address_in = 16#08C9# else
		x"059D" when address_in = 16#08CA# else
		x"F300" when address_in = 16#08CB# else
		x"2DBF" when address_in = 16#08CC# else
		x"2DAE" when address_in = 16#08CD# else
		x"918D" when address_in = 16#08CE# else
		x"919C" when address_in = 16#08CF# else
		x"158C" when address_in = 16#08D0# else
		x"059D" when address_in = 16#08D1# else
		x"F458" when address_in = 16#08D2# else
		x"2DFF" when address_in = 16#08D3# else
		x"2DEE" when address_in = 16#08D4# else
		x"80E5" when address_in = 16#08D5# else
		x"80F6" when address_in = 16#08D6# else
		x"9180" when address_in = 16#08D7# else
		x"007C" when address_in = 16#08D8# else
		x"9190" when address_in = 16#08D9# else
		x"007D" when address_in = 16#08DA# else
		x"16E8" when address_in = 16#08DB# else
		x"06F9" when address_in = 16#08DC# else
		x"F671" when address_in = 16#08DD# else
		x"9180" when address_in = 16#08DE# else
		x"007C" when address_in = 16#08DF# else
		x"9190" when address_in = 16#08E0# else
		x"007D" when address_in = 16#08E1# else
		x"16E8" when address_in = 16#08E2# else
		x"06F9" when address_in = 16#08E3# else
		x"F421" when address_in = 16#08E4# else
		x"BF0F" when address_in = 16#08E5# else
		x"E080" when address_in = 16#08E6# else
		x"E090" when address_in = 16#08E7# else
		x"C04F" when address_in = 16#08E8# else
		x"2DBF" when address_in = 16#08E9# else
		x"2DAE" when address_in = 16#08EA# else
		x"918D" when address_in = 16#08EB# else
		x"919C" when address_in = 16#08EC# else
		x"9711" when address_in = 16#08ED# else
		x"16C8" when address_in = 16#08EE# else
		x"06D9" when address_in = 16#08EF# else
		x"F498" when address_in = 16#08F0# else
		x"2DFD" when address_in = 16#08F1# else
		x"2DEC" when address_in = 16#08F2# else
		x"E0C3" when address_in = 16#08F3# else
		x"0FEE" when address_in = 16#08F4# else
		x"1FFF" when address_in = 16#08F5# else
		x"95CA" when address_in = 16#08F6# else
		x"F7E1" when address_in = 16#08F7# else
		x"0DEE" when address_in = 16#08F8# else
		x"1DFF" when address_in = 16#08F9# else
		x"198C" when address_in = 16#08FA# else
		x"099D" when address_in = 16#08FB# else
		x"8391" when address_in = 16#08FC# else
		x"8380" when address_in = 16#08FD# else
		x"92CD" when address_in = 16#08FE# else
		x"92DC" when address_in = 16#08FF# else
		x"2F8E" when address_in = 16#0900# else
		x"2F9F" when address_in = 16#0901# else
		x"940E" when address_in = 16#0902# else
		x"07D3" when address_in = 16#0903# else
		x"2D9F" when address_in = 16#0904# else
		x"2D8E" when address_in = 16#0905# else
		x"940E" when address_in = 16#0906# else
		x"062C" when address_in = 16#0907# else
		x"2DFF" when address_in = 16#0908# else
		x"2DEE" when address_in = 16#0909# else
		x"8180" when address_in = 16#090A# else
		x"8191" when address_in = 16#090B# else
		x"6890" when address_in = 16#090C# else
		x"8391" when address_in = 16#090D# else
		x"8380" when address_in = 16#090E# else
		x"82B2" when address_in = 16#090F# else
		x"3017" when address_in = 16#0910# else
		x"F429" when address_in = 16#0911# else
		x"2D8B" when address_in = 16#0912# else
		x"940E" when address_in = 16#0913# else
		x"2D9E" when address_in = 16#0914# else
		x"2F48" when address_in = 16#0915# else
		x"C001" when address_in = 16#0916# else
		x"2F41" when address_in = 16#0917# else
		x"2F14" when address_in = 16#0918# else
		x"7017" when address_in = 16#0919# else
		x"2F81" when address_in = 16#091A# else
		x"6088" when address_in = 16#091B# else
		x"2F48" when address_in = 16#091C# else
		x"E068" when address_in = 16#091D# else
		x"E070" when address_in = 16#091E# else
		x"2D9F" when address_in = 16#091F# else
		x"2D8E" when address_in = 16#0920# else
		x"940E" when address_in = 16#0921# else
		x"0A4B" when address_in = 16#0922# else
		x"E0F3" when address_in = 16#0923# else
		x"0CCC" when address_in = 16#0924# else
		x"1CDD" when address_in = 16#0925# else
		x"95FA" when address_in = 16#0926# else
		x"F7E1" when address_in = 16#0927# else
		x"EF88" when address_in = 16#0928# else
		x"EF9F" when address_in = 16#0929# else
		x"0EC8" when address_in = 16#092A# else
		x"1ED9" when address_in = 16#092B# else
		x"2F41" when address_in = 16#092C# else
		x"2D7D" when address_in = 16#092D# else
		x"2D6C" when address_in = 16#092E# else
		x"2D9F" when address_in = 16#092F# else
		x"2D8E" when address_in = 16#0930# else
		x"9608" when address_in = 16#0931# else
		x"940E" when address_in = 16#0932# else
		x"0A4B" when address_in = 16#0933# else
		x"BF0F" when address_in = 16#0934# else
		x"2D9F" when address_in = 16#0935# else
		x"2D8E" when address_in = 16#0936# else
		x"9603" when address_in = 16#0937# else
		x"91DF" when address_in = 16#0938# else
		x"91CF" when address_in = 16#0939# else
		x"911F" when address_in = 16#093A# else
		x"910F" when address_in = 16#093B# else
		x"90FF" when address_in = 16#093C# else
		x"90EF" when address_in = 16#093D# else
		x"90DF" when address_in = 16#093E# else
		x"90CF" when address_in = 16#093F# else
		x"90BF" when address_in = 16#0940# else
		x"9508" when address_in = 16#0941# else
		x"930F" when address_in = 16#0942# else
		x"931F" when address_in = 16#0943# else
		x"93CF" when address_in = 16#0944# else
		x"93DF" when address_in = 16#0945# else
		x"2F08" when address_in = 16#0946# else
		x"E9C0" when address_in = 16#0947# else
		x"E0D1" when address_in = 16#0948# else
		x"B71F" when address_in = 16#0949# else
		x"94F8" when address_in = 16#094A# else
		x"9180" when address_in = 16#094B# else
		x"007C" when address_in = 16#094C# else
		x"9190" when address_in = 16#094D# else
		x"007D" when address_in = 16#094E# else
		x"17C8" when address_in = 16#094F# else
		x"07D9" when address_in = 16#0950# else
		x"F0F9" when address_in = 16#0951# else
		x"8188" when address_in = 16#0952# else
		x"8199" when address_in = 16#0953# else
		x"FF97" when address_in = 16#0954# else
		x"C011" when address_in = 16#0955# else
		x"818A" when address_in = 16#0956# else
		x"1780" when address_in = 16#0957# else
		x"F471" when address_in = 16#0958# else
		x"B184" when address_in = 16#0959# else
		x"2799" when address_in = 16#095A# else
		x"718E" when address_in = 16#095B# else
		x"7090" when address_in = 16#095C# else
		x"9595" when address_in = 16#095D# else
		x"9587" when address_in = 16#095E# else
		x"9595" when address_in = 16#095F# else
		x"9587" when address_in = 16#0960# else
		x"2F68" when address_in = 16#0961# else
		x"2F8C" when address_in = 16#0962# else
		x"2F9D" when address_in = 16#0963# else
		x"9603" when address_in = 16#0964# else
		x"940E" when address_in = 16#0965# else
		x"07EC" when address_in = 16#0966# else
		x"8188" when address_in = 16#0967# else
		x"8199" when address_in = 16#0968# else
		x"E033" when address_in = 16#0969# else
		x"0F88" when address_in = 16#096A# else
		x"1F99" when address_in = 16#096B# else
		x"953A" when address_in = 16#096C# else
		x"F7E1" when address_in = 16#096D# else
		x"0FC8" when address_in = 16#096E# else
		x"1FD9" when address_in = 16#096F# else
		x"CFDA" when address_in = 16#0970# else
		x"BF1F" when address_in = 16#0971# else
		x"E080" when address_in = 16#0972# else
		x"E090" when address_in = 16#0973# else
		x"91DF" when address_in = 16#0974# else
		x"91CF" when address_in = 16#0975# else
		x"911F" when address_in = 16#0976# else
		x"910F" when address_in = 16#0977# else
		x"9508" when address_in = 16#0978# else
		x"92EF" when address_in = 16#0979# else
		x"92FF" when address_in = 16#097A# else
		x"930F" when address_in = 16#097B# else
		x"931F" when address_in = 16#097C# else
		x"E900" when address_in = 16#097D# else
		x"E011" when address_in = 16#097E# else
		x"2CE1" when address_in = 16#097F# else
		x"E0F8" when address_in = 16#0980# else
		x"2EFF" when address_in = 16#0981# else
		x"0EE0" when address_in = 16#0982# else
		x"1EF1" when address_in = 16#0983# else
		x"9310" when address_in = 16#0984# else
		x"007B" when address_in = 16#0985# else
		x"9300" when address_in = 16#0986# else
		x"007A" when address_in = 16#0987# else
		x"EF4F" when address_in = 16#0988# else
		x"E050" when address_in = 16#0989# else
		x"9350" when address_in = 16#098A# else
		x"007F" when address_in = 16#098B# else
		x"9340" when address_in = 16#098C# else
		x"007E" when address_in = 16#098D# else
		x"2F31" when address_in = 16#098E# else
		x"2F20" when address_in = 16#098F# else
		x"5028" when address_in = 16#0990# else
		x"4F38" when address_in = 16#0991# else
		x"9330" when address_in = 16#0992# else
		x"007D" when address_in = 16#0993# else
		x"9320" when address_in = 16#0994# else
		x"007C" when address_in = 16#0995# else
		x"E080" when address_in = 16#0996# else
		x"E890" when address_in = 16#0997# else
		x"9390" when address_in = 16#0998# else
		x"0989" when address_in = 16#0999# else
		x"9380" when address_in = 16#099A# else
		x"0988" when address_in = 16#099B# else
		x"9330" when address_in = 16#099C# else
		x"098C" when address_in = 16#099D# else
		x"9320" when address_in = 16#099E# else
		x"098B" when address_in = 16#099F# else
		x"9330" when address_in = 16#09A0# else
		x"098E" when address_in = 16#09A1# else
		x"9320" when address_in = 16#09A2# else
		x"098D" when address_in = 16#09A3# else
		x"9350" when address_in = 16#09A4# else
		x"0191" when address_in = 16#09A5# else
		x"9340" when address_in = 16#09A6# else
		x"0190" when address_in = 16#09A7# else
		x"2F91" when address_in = 16#09A8# else
		x"2F80" when address_in = 16#09A9# else
		x"940E" when address_in = 16#09AA# else
		x"07D3" when address_in = 16#09AB# else
		x"940E" when address_in = 16#09AC# else
		x"0A41" when address_in = 16#09AD# else
		x"9180" when address_in = 16#09AE# else
		x"007E" when address_in = 16#09AF# else
		x"9190" when address_in = 16#09B0# else
		x"007F" when address_in = 16#09B1# else
		x"E0E3" when address_in = 16#09B2# else
		x"0F88" when address_in = 16#09B3# else
		x"1F99" when address_in = 16#09B4# else
		x"95EA" when address_in = 16#09B5# else
		x"F7E1" when address_in = 16#09B6# else
		x"E04F" when address_in = 16#09B7# else
		x"2F68" when address_in = 16#09B8# else
		x"2F79" when address_in = 16#09B9# else
		x"9180" when address_in = 16#09BA# else
		x"007A" when address_in = 16#09BB# else
		x"9190" when address_in = 16#09BC# else
		x"007B" when address_in = 16#09BD# else
		x"940E" when address_in = 16#09BE# else
		x"0A4B" when address_in = 16#09BF# else
		x"9310" when address_in = 16#09C0# else
		x"0172" when address_in = 16#09C1# else
		x"9300" when address_in = 16#09C2# else
		x"0171" when address_in = 16#09C3# else
		x"B184" when address_in = 16#09C4# else
		x"718F" when address_in = 16#09C5# else
		x"B984" when address_in = 16#09C6# else
		x"B184" when address_in = 16#09C7# else
		x"6680" when address_in = 16#09C8# else
		x"B984" when address_in = 16#09C9# else
		x"9821" when address_in = 16#09CA# else
		x"B908" when address_in = 16#09CB# else
		x"2F81" when address_in = 16#09CC# else
		x"2799" when address_in = 16#09CD# else
		x"B987" when address_in = 16#09CE# else
		x"B8E6" when address_in = 16#09CF# else
		x"2D8F" when address_in = 16#09D0# else
		x"2799" when address_in = 16#09D1# else
		x"B985" when address_in = 16#09D2# else
		x"E980" when address_in = 16#09D3# else
		x"E099" when address_in = 16#09D4# else
		x"BB8D" when address_in = 16#09D5# else
		x"2F89" when address_in = 16#09D6# else
		x"2799" when address_in = 16#09D7# else
		x"BB8E" when address_in = 16#09D8# else
		x"9A20" when address_in = 16#09D9# else
		x"911F" when address_in = 16#09DA# else
		x"910F" when address_in = 16#09DB# else
		x"90FF" when address_in = 16#09DC# else
		x"90EF" when address_in = 16#09DD# else
		x"9508" when address_in = 16#09DE# else
		x"93CF" when address_in = 16#09DF# else
		x"93DF" when address_in = 16#09E0# else
		x"E081" when address_in = 16#09E1# else
		x"940E" when address_in = 16#09E2# else
		x"26CF" when address_in = 16#09E3# else
		x"E082" when address_in = 16#09E4# else
		x"940E" when address_in = 16#09E5# else
		x"26CF" when address_in = 16#09E6# else
		x"E083" when address_in = 16#09E7# else
		x"940E" when address_in = 16#09E8# else
		x"26CF" when address_in = 16#09E9# else
		x"EFCF" when address_in = 16#09EA# else
		x"EFDF" when address_in = 16#09EB# else
		x"95A8" when address_in = 16#09EC# else
		x"9720" when address_in = 16#09ED# else
		x"F449" when address_in = 16#09EE# else
		x"E087" when address_in = 16#09EF# else
		x"940E" when address_in = 16#09F0# else
		x"26CF" when address_in = 16#09F1# else
		x"E088" when address_in = 16#09F2# else
		x"940E" when address_in = 16#09F3# else
		x"26CF" when address_in = 16#09F4# else
		x"E089" when address_in = 16#09F5# else
		x"940E" when address_in = 16#09F6# else
		x"26CF" when address_in = 16#09F7# else
		x"9721" when address_in = 16#09F8# else
		x"CFF2" when address_in = 16#09F9# else
		x"940E" when address_in = 16#09FA# else
		x"09DF" when address_in = 16#09FB# else
		x"2799" when address_in = 16#09FC# else
		x"FD87" when address_in = 16#09FD# else
		x"9590" when address_in = 16#09FE# else
		x"9508" when address_in = 16#09FF# else
		x"92EF" when address_in = 16#0A00# else
		x"92FF" when address_in = 16#0A01# else
		x"930F" when address_in = 16#0A02# else
		x"931F" when address_in = 16#0A03# else
		x"93CF" when address_in = 16#0A04# else
		x"93DF" when address_in = 16#0A05# else
		x"2F08" when address_in = 16#0A06# else
		x"2F19" when address_in = 16#0A07# else
		x"2EF6" when address_in = 16#0A08# else
		x"940E" when address_in = 16#0A09# else
		x"0B5D" when address_in = 16#0A0A# else
		x"2EE8" when address_in = 16#0A0B# else
		x"2D4F" when address_in = 16#0A0C# else
		x"2F68" when address_in = 16#0A0D# else
		x"2F91" when address_in = 16#0A0E# else
		x"2F80" when address_in = 16#0A0F# else
		x"940E" when address_in = 16#0A10# else
		x"0889" when address_in = 16#0A11# else
		x"2FD9" when address_in = 16#0A12# else
		x"2FC8" when address_in = 16#0A13# else
		x"2B89" when address_in = 16#0A14# else
		x"F419" when address_in = 16#0A15# else
		x"2D8E" when address_in = 16#0A16# else
		x"940E" when address_in = 16#0A17# else
		x"09FA" when address_in = 16#0A18# else
		x"2F8C" when address_in = 16#0A19# else
		x"2F9D" when address_in = 16#0A1A# else
		x"91DF" when address_in = 16#0A1B# else
		x"91CF" when address_in = 16#0A1C# else
		x"911F" when address_in = 16#0A1D# else
		x"910F" when address_in = 16#0A1E# else
		x"90FF" when address_in = 16#0A1F# else
		x"90EF" when address_in = 16#0A20# else
		x"9508" when address_in = 16#0A21# else
		x"940E" when address_in = 16#0A22# else
		x"07EC" when address_in = 16#0A23# else
		x"9508" when address_in = 16#0A24# else
		x"92FF" when address_in = 16#0A25# else
		x"930F" when address_in = 16#0A26# else
		x"931F" when address_in = 16#0A27# else
		x"93CF" when address_in = 16#0A28# else
		x"2F08" when address_in = 16#0A29# else
		x"2F19" when address_in = 16#0A2A# else
		x"2EF6" when address_in = 16#0A2B# else
		x"940E" when address_in = 16#0A2C# else
		x"0B5D" when address_in = 16#0A2D# else
		x"2FC8" when address_in = 16#0A2E# else
		x"2D4F" when address_in = 16#0A2F# else
		x"2F68" when address_in = 16#0A30# else
		x"2F91" when address_in = 16#0A31# else
		x"2F80" when address_in = 16#0A32# else
		x"940E" when address_in = 16#0A33# else
		x"0700" when address_in = 16#0A34# else
		x"2388" when address_in = 16#0A35# else
		x"F019" when address_in = 16#0A36# else
		x"2F8C" when address_in = 16#0A37# else
		x"940E" when address_in = 16#0A38# else
		x"09FA" when address_in = 16#0A39# else
		x"E080" when address_in = 16#0A3A# else
		x"E090" when address_in = 16#0A3B# else
		x"91CF" when address_in = 16#0A3C# else
		x"911F" when address_in = 16#0A3D# else
		x"910F" when address_in = 16#0A3E# else
		x"90FF" when address_in = 16#0A3F# else
		x"9508" when address_in = 16#0A40# else
		x"EF8F" when address_in = 16#0A41# else
		x"E9E0" when address_in = 16#0A42# else
		x"E0F9" when address_in = 16#0A43# else
		x"9381" when address_in = 16#0A44# else
		x"E09A" when address_in = 16#0A45# else
		x"38EF" when address_in = 16#0A46# else
		x"07F9" when address_in = 16#0A47# else
		x"F3D9" when address_in = 16#0A48# else
		x"F3D0" when address_in = 16#0A49# else
		x"9508" when address_in = 16#0A4A# else
		x"93CF" when address_in = 16#0A4B# else
		x"2F28" when address_in = 16#0A4C# else
		x"2F39" when address_in = 16#0A4D# else
		x"2FC4" when address_in = 16#0A4E# else
		x"1561" when address_in = 16#0A4F# else
		x"0571" when address_in = 16#0A50# else
		x"F409" when address_in = 16#0A51# else
		x"C04B" when address_in = 16#0A52# else
		x"2F97" when address_in = 16#0A53# else
		x"2F86" when address_in = 16#0A54# else
		x"7087" when address_in = 16#0A55# else
		x"7F98" when address_in = 16#0A56# else
		x"2B89" when address_in = 16#0A57# else
		x"F009" when address_in = 16#0A58# else
		x"C044" when address_in = 16#0A59# else
		x"E043" when address_in = 16#0A5A# else
		x"9576" when address_in = 16#0A5B# else
		x"9567" when address_in = 16#0A5C# else
		x"954A" when address_in = 16#0A5D# else
		x"F7E1" when address_in = 16#0A5E# else
		x"9180" when address_in = 16#0A5F# else
		x"0171" when address_in = 16#0A60# else
		x"9190" when address_in = 16#0A61# else
		x"0172" when address_in = 16#0A62# else
		x"1B28" when address_in = 16#0A63# else
		x"0B39" when address_in = 16#0A64# else
		x"2FB3" when address_in = 16#0A65# else
		x"2FA2" when address_in = 16#0A66# else
		x"E094" when address_in = 16#0A67# else
		x"95B6" when address_in = 16#0A68# else
		x"95A7" when address_in = 16#0A69# else
		x"959A" when address_in = 16#0A6A# else
		x"F7E1" when address_in = 16#0A6B# else
		x"9536" when address_in = 16#0A6C# else
		x"9527" when address_in = 16#0A6D# else
		x"2FFB" when address_in = 16#0A6E# else
		x"2FEA" when address_in = 16#0A6F# else
		x"57E0" when address_in = 16#0A70# else
		x"4FF6" when address_in = 16#0A71# else
		x"8150" when address_in = 16#0A72# else
		x"7024" when address_in = 16#0A73# else
		x"7030" when address_in = 16#0A74# else
		x"E08F" when address_in = 16#0A75# else
		x"E090" when address_in = 16#0A76# else
		x"2E02" when address_in = 16#0A77# else
		x"C002" when address_in = 16#0A78# else
		x"0F88" when address_in = 16#0A79# else
		x"1F99" when address_in = 16#0A7A# else
		x"940A" when address_in = 16#0A7B# else
		x"F7E2" when address_in = 16#0A7C# else
		x"2F48" when address_in = 16#0A7D# else
		x"2F8C" when address_in = 16#0A7E# else
		x"2799" when address_in = 16#0A7F# else
		x"C002" when address_in = 16#0A80# else
		x"0F88" when address_in = 16#0A81# else
		x"1F99" when address_in = 16#0A82# else
		x"952A" when address_in = 16#0A83# else
		x"F7E2" when address_in = 16#0A84# else
		x"2F98" when address_in = 16#0A85# else
		x"1561" when address_in = 16#0A86# else
		x"0571" when address_in = 16#0A87# else
		x"F091" when address_in = 16#0A88# else
		x"2F84" when address_in = 16#0A89# else
		x"9580" when address_in = 16#0A8A# else
		x"2358" when address_in = 16#0A8B# else
		x"2B59" when address_in = 16#0A8C# else
		x"5061" when address_in = 16#0A8D# else
		x"4070" when address_in = 16#0A8E# else
		x"9542" when address_in = 16#0A8F# else
		x"7F40" when address_in = 16#0A90# else
		x"9592" when address_in = 16#0A91# else
		x"7F90" when address_in = 16#0A92# else
		x"2344" when address_in = 16#0A93# else
		x"F789" when address_in = 16#0A94# else
		x"9351" when address_in = 16#0A95# else
		x"9611" when address_in = 16#0A96# else
		x"8150" when address_in = 16#0A97# else
		x"E04F" when address_in = 16#0A98# else
		x"2F9C" when address_in = 16#0A99# else
		x"CFEB" when address_in = 16#0A9A# else
		x"57A0" when address_in = 16#0A9B# else
		x"4FB6" when address_in = 16#0A9C# else
		x"935C" when address_in = 16#0A9D# else
		x"91CF" when address_in = 16#0A9E# else
		x"9508" when address_in = 16#0A9F# else
		x"92FF" when address_in = 16#0AA0# else
		x"930F" when address_in = 16#0AA1# else
		x"931F" when address_in = 16#0AA2# else
		x"93CF" when address_in = 16#0AA3# else
		x"93DF" when address_in = 16#0AA4# else
		x"2EF6" when address_in = 16#0AA5# else
		x"2F04" when address_in = 16#0AA6# else
		x"2F12" when address_in = 16#0AA7# else
		x"E0C0" when address_in = 16#0AA8# else
		x"E0D0" when address_in = 16#0AA9# else
		x"9120" when address_in = 16#0AAA# else
		x"0171" when address_in = 16#0AAB# else
		x"9130" when address_in = 16#0AAC# else
		x"0172" when address_in = 16#0AAD# else
		x"1B82" when address_in = 16#0AAE# else
		x"0B93" when address_in = 16#0AAF# else
		x"2FB9" when address_in = 16#0AB0# else
		x"2FA8" when address_in = 16#0AB1# else
		x"E064" when address_in = 16#0AB2# else
		x"95B6" when address_in = 16#0AB3# else
		x"95A7" when address_in = 16#0AB4# else
		x"956A" when address_in = 16#0AB5# else
		x"F7E1" when address_in = 16#0AB6# else
		x"2F28" when address_in = 16#0AB7# else
		x"2F39" when address_in = 16#0AB8# else
		x"9536" when address_in = 16#0AB9# else
		x"9527" when address_in = 16#0ABA# else
		x"2FFB" when address_in = 16#0ABB# else
		x"2FEA" when address_in = 16#0ABC# else
		x"57E0" when address_in = 16#0ABD# else
		x"4FF6" when address_in = 16#0ABE# else
		x"8150" when address_in = 16#0ABF# else
		x"2D8F" when address_in = 16#0AC0# else
		x"2799" when address_in = 16#0AC1# else
		x"7024" when address_in = 16#0AC2# else
		x"7030" when address_in = 16#0AC3# else
		x"2E02" when address_in = 16#0AC4# else
		x"C002" when address_in = 16#0AC5# else
		x"0F88" when address_in = 16#0AC6# else
		x"1F99" when address_in = 16#0AC7# else
		x"940A" when address_in = 16#0AC8# else
		x"F7E2" when address_in = 16#0AC9# else
		x"2F68" when address_in = 16#0ACA# else
		x"2F84" when address_in = 16#0ACB# else
		x"2799" when address_in = 16#0ACC# else
		x"2E02" when address_in = 16#0ACD# else
		x"C002" when address_in = 16#0ACE# else
		x"0F88" when address_in = 16#0ACF# else
		x"1F99" when address_in = 16#0AD0# else
		x"940A" when address_in = 16#0AD1# else
		x"F7E2" when address_in = 16#0AD2# else
		x"2F78" when address_in = 16#0AD3# else
		x"2F81" when address_in = 16#0AD4# else
		x"2799" when address_in = 16#0AD5# else
		x"2E02" when address_in = 16#0AD6# else
		x"C002" when address_in = 16#0AD7# else
		x"0F88" when address_in = 16#0AD8# else
		x"1F99" when address_in = 16#0AD9# else
		x"940A" when address_in = 16#0ADA# else
		x"F7E2" when address_in = 16#0ADB# else
		x"2F48" when address_in = 16#0ADC# else
		x"E08F" when address_in = 16#0ADD# else
		x"E090" when address_in = 16#0ADE# else
		x"C002" when address_in = 16#0ADF# else
		x"0F88" when address_in = 16#0AE0# else
		x"1F99" when address_in = 16#0AE1# else
		x"952A" when address_in = 16#0AE2# else
		x"F7E2" when address_in = 16#0AE3# else
		x"2F98" when address_in = 16#0AE4# else
		x"2F85" when address_in = 16#0AE5# else
		x"2386" when address_in = 16#0AE6# else
		x"1787" when address_in = 16#0AE7# else
		x"F4B1" when address_in = 16#0AE8# else
		x"2F89" when address_in = 16#0AE9# else
		x"9580" when address_in = 16#0AEA# else
		x"2358" when address_in = 16#0AEB# else
		x"2B54" when address_in = 16#0AEC# else
		x"9621" when address_in = 16#0AED# else
		x"9562" when address_in = 16#0AEE# else
		x"7F60" when address_in = 16#0AEF# else
		x"9572" when address_in = 16#0AF0# else
		x"7F70" when address_in = 16#0AF1# else
		x"9542" when address_in = 16#0AF2# else
		x"7F40" when address_in = 16#0AF3# else
		x"9592" when address_in = 16#0AF4# else
		x"7F90" when address_in = 16#0AF5# else
		x"F771" when address_in = 16#0AF6# else
		x"9351" when address_in = 16#0AF7# else
		x"9611" when address_in = 16#0AF8# else
		x"8150" when address_in = 16#0AF9# else
		x"2D6F" when address_in = 16#0AFA# else
		x"2F70" when address_in = 16#0AFB# else
		x"2F41" when address_in = 16#0AFC# else
		x"E09F" when address_in = 16#0AFD# else
		x"CFE6" when address_in = 16#0AFE# else
		x"57A0" when address_in = 16#0AFF# else
		x"4FB6" when address_in = 16#0B00# else
		x"935C" when address_in = 16#0B01# else
		x"2F8C" when address_in = 16#0B02# else
		x"2F9D" when address_in = 16#0B03# else
		x"91DF" when address_in = 16#0B04# else
		x"91CF" when address_in = 16#0B05# else
		x"911F" when address_in = 16#0B06# else
		x"910F" when address_in = 16#0B07# else
		x"90FF" when address_in = 16#0B08# else
		x"9508" when address_in = 16#0B09# else
		x"940E" when address_in = 16#0B0A# else
		x"0621" when address_in = 16#0B0B# else
		x"940E" when address_in = 16#0B0C# else
		x"0D10" when address_in = 16#0B0D# else
		x"9508" when address_in = 16#0B0E# else
		x"2FF7" when address_in = 16#0B0F# else
		x"2FE6" when address_in = 16#0B10# else
		x"8186" when address_in = 16#0B11# else
		x"2388" when address_in = 16#0B12# else
		x"F419" when address_in = 16#0B13# else
		x"E080" when address_in = 16#0B14# else
		x"E090" when address_in = 16#0B15# else
		x"9508" when address_in = 16#0B16# else
		x"EE8A" when address_in = 16#0B17# else
		x"EF9F" when address_in = 16#0B18# else
		x"9508" when address_in = 16#0B19# else
		x"3084" when address_in = 16#0B1A# else
		x"F458" when address_in = 16#0B1B# else
		x"2FE8" when address_in = 16#0B1C# else
		x"27FF" when address_in = 16#0B1D# else
		x"0FEE" when address_in = 16#0B1E# else
		x"1FFF" when address_in = 16#0B1F# else
		x"56E7" when address_in = 16#0B20# else
		x"4FFF" when address_in = 16#0B21# else
		x"8371" when address_in = 16#0B22# else
		x"8360" when address_in = 16#0B23# else
		x"E081" when address_in = 16#0B24# else
		x"9380" when address_in = 16#0B25# else
		x"0080" when address_in = 16#0B26# else
		x"9508" when address_in = 16#0B27# else
		x"2F98" when address_in = 16#0B28# else
		x"7083" when address_in = 16#0B29# else
		x"2FE8" when address_in = 16#0B2A# else
		x"27FF" when address_in = 16#0B2B# else
		x"0FEE" when address_in = 16#0B2C# else
		x"1FFF" when address_in = 16#0B2D# else
		x"57EA" when address_in = 16#0B2E# else
		x"4FFE" when address_in = 16#0B2F# else
		x"9001" when address_in = 16#0B30# else
		x"81F0" when address_in = 16#0B31# else
		x"2DE0" when address_in = 16#0B32# else
		x"9730" when address_in = 16#0B33# else
		x"F031" when address_in = 16#0B34# else
		x"8184" when address_in = 16#0B35# else
		x"1789" when address_in = 16#0B36# else
		x"F7C1" when address_in = 16#0B37# else
		x"2F8E" when address_in = 16#0B38# else
		x"2F9F" when address_in = 16#0B39# else
		x"9508" when address_in = 16#0B3A# else
		x"E080" when address_in = 16#0B3B# else
		x"E090" when address_in = 16#0B3C# else
		x"9508" when address_in = 16#0B3D# else
		x"940E" when address_in = 16#0B3E# else
		x"0B28" when address_in = 16#0B3F# else
		x"2FF9" when address_in = 16#0B40# else
		x"2FE8" when address_in = 16#0B41# else
		x"9700" when address_in = 16#0B42# else
		x"F409" when address_in = 16#0B43# else
		x"9508" when address_in = 16#0B44# else
		x"8186" when address_in = 16#0B45# else
		x"8197" when address_in = 16#0B46# else
		x"9508" when address_in = 16#0B47# else
		x"9180" when address_in = 16#0B48# else
		x"0173" when address_in = 16#0B49# else
		x"940E" when address_in = 16#0B4A# else
		x"0B28" when address_in = 16#0B4B# else
		x"2FF9" when address_in = 16#0B4C# else
		x"2FE8" when address_in = 16#0B4D# else
		x"9700" when address_in = 16#0B4E# else
		x"F409" when address_in = 16#0B4F# else
		x"9508" when address_in = 16#0B50# else
		x"8186" when address_in = 16#0B51# else
		x"8197" when address_in = 16#0B52# else
		x"9508" when address_in = 16#0B53# else
		x"9190" when address_in = 16#0B54# else
		x"0173" when address_in = 16#0B55# else
		x"3F8F" when address_in = 16#0B56# else
		x"F011" when address_in = 16#0B57# else
		x"9380" when address_in = 16#0B58# else
		x"0173" when address_in = 16#0B59# else
		x"2F89" when address_in = 16#0B5A# else
		x"2799" when address_in = 16#0B5B# else
		x"9508" when address_in = 16#0B5C# else
		x"9180" when address_in = 16#0B5D# else
		x"0173" when address_in = 16#0B5E# else
		x"2799" when address_in = 16#0B5F# else
		x"9508" when address_in = 16#0B60# else
		x"E886" when address_in = 16#0B61# else
		x"E091" when address_in = 16#0B62# else
		x"9508" when address_in = 16#0B63# else
		x"92CF" when address_in = 16#0B64# else
		x"92DF" when address_in = 16#0B65# else
		x"92EF" when address_in = 16#0B66# else
		x"92FF" when address_in = 16#0B67# else
		x"930F" when address_in = 16#0B68# else
		x"931F" when address_in = 16#0B69# else
		x"93CF" when address_in = 16#0B6A# else
		x"93DF" when address_in = 16#0B6B# else
		x"2FD9" when address_in = 16#0B6C# else
		x"2FC8" when address_in = 16#0B6D# else
		x"2EE6" when address_in = 16#0B6E# else
		x"2EF7" when address_in = 16#0B6F# else
		x"2F04" when address_in = 16#0B70# else
		x"2F15" when address_in = 16#0B71# else
		x"2EC2" when address_in = 16#0B72# else
		x"818C" when address_in = 16#0B73# else
		x"E033" when address_in = 16#0B74# else
		x"2ED3" when address_in = 16#0B75# else
		x"22D8" when address_in = 16#0B76# else
		x"940E" when address_in = 16#0B77# else
		x"0B28" when address_in = 16#0B78# else
		x"2B89" when address_in = 16#0B79# else
		x"F019" when address_in = 16#0B7A# else
		x"EE8F" when address_in = 16#0B7B# else
		x"EF9F" when address_in = 16#0B7C# else
		x"C03D" when address_in = 16#0B7D# else
		x"2D8E" when address_in = 16#0B7E# else
		x"2D9F" when address_in = 16#0B7F# else
		x"27AA" when address_in = 16#0B80# else
		x"27BB" when address_in = 16#0B81# else
		x"0F88" when address_in = 16#0B82# else
		x"1F99" when address_in = 16#0B83# else
		x"1FAA" when address_in = 16#0B84# else
		x"1FBB" when address_in = 16#0B85# else
		x"9602" when address_in = 16#0B86# else
		x"1DA1" when address_in = 16#0B87# else
		x"1DB1" when address_in = 16#0B88# else
		x"BFAB" when address_in = 16#0B89# else
		x"2FF9" when address_in = 16#0B8A# else
		x"2FE8" when address_in = 16#0B8B# else
		x"95D8" when address_in = 16#0B8C# else
		x"2D60" when address_in = 16#0B8D# else
		x"2366" when address_in = 16#0B8E# else
		x"F029" when address_in = 16#0B8F# else
		x"818C" when address_in = 16#0B90# else
		x"940E" when address_in = 16#0B91# else
		x"1C51" when address_in = 16#0B92# else
		x"2388" when address_in = 16#0B93# else
		x"F10C" when address_in = 16#0B94# else
		x"2F8C" when address_in = 16#0B95# else
		x"2F9D" when address_in = 16#0B96# else
		x"940E" when address_in = 16#0B97# else
		x"1A0E" when address_in = 16#0B98# else
		x"B78F" when address_in = 16#0B99# else
		x"94F8" when address_in = 16#0B9A# else
		x"2DED" when address_in = 16#0B9B# else
		x"27FF" when address_in = 16#0B9C# else
		x"0FEE" when address_in = 16#0B9D# else
		x"1FFF" when address_in = 16#0B9E# else
		x"57EA" when address_in = 16#0B9F# else
		x"4FFE" when address_in = 16#0BA0# else
		x"8120" when address_in = 16#0BA1# else
		x"8131" when address_in = 16#0BA2# else
		x"8339" when address_in = 16#0BA3# else
		x"8328" when address_in = 16#0BA4# else
		x"83D1" when address_in = 16#0BA5# else
		x"83C0" when address_in = 16#0BA6# else
		x"BF8F" when address_in = 16#0BA7# else
		x"E884" when address_in = 16#0BA8# else
		x"2EE8" when address_in = 16#0BA9# else
		x"2CF1" when address_in = 16#0BAA# else
		x"2D2C" when address_in = 16#0BAB# else
		x"E040" when address_in = 16#0BAC# else
		x"E062" when address_in = 16#0BAD# else
		x"818C" when address_in = 16#0BAE# else
		x"940E" when address_in = 16#0BAF# else
		x"105C" when address_in = 16#0BB0# else
		x"2388" when address_in = 16#0BB1# else
		x"F031" when address_in = 16#0BB2# else
		x"818C" when address_in = 16#0BB3# else
		x"940E" when address_in = 16#0BB4# else
		x"1BAF" when address_in = 16#0BB5# else
		x"EF84" when address_in = 16#0BB6# else
		x"EF9F" when address_in = 16#0BB7# else
		x"C002" when address_in = 16#0BB8# else
		x"E080" when address_in = 16#0BB9# else
		x"E090" when address_in = 16#0BBA# else
		x"91DF" when address_in = 16#0BBB# else
		x"91CF" when address_in = 16#0BBC# else
		x"911F" when address_in = 16#0BBD# else
		x"910F" when address_in = 16#0BBE# else
		x"90FF" when address_in = 16#0BBF# else
		x"90EF" when address_in = 16#0BC0# else
		x"90DF" when address_in = 16#0BC1# else
		x"90CF" when address_in = 16#0BC2# else
		x"9508" when address_in = 16#0BC3# else
		x"93CF" when address_in = 16#0BC4# else
		x"93DF" when address_in = 16#0BC5# else
		x"2FD9" when address_in = 16#0BC6# else
		x"2FC8" when address_in = 16#0BC7# else
		x"1561" when address_in = 16#0BC8# else
		x"0571" when address_in = 16#0BC9# else
		x"F079" when address_in = 16#0BCA# else
		x"2F86" when address_in = 16#0BCB# else
		x"2F97" when address_in = 16#0BCC# else
		x"27AA" when address_in = 16#0BCD# else
		x"27BB" when address_in = 16#0BCE# else
		x"0F88" when address_in = 16#0BCF# else
		x"1F99" when address_in = 16#0BD0# else
		x"1FAA" when address_in = 16#0BD1# else
		x"1FBB" when address_in = 16#0BD2# else
		x"BFAB" when address_in = 16#0BD3# else
		x"2FF9" when address_in = 16#0BD4# else
		x"2FE8" when address_in = 16#0BD5# else
		x"95D8" when address_in = 16#0BD6# else
		x"2D80" when address_in = 16#0BD7# else
		x"3E80" when address_in = 16#0BD8# else
		x"F018" when address_in = 16#0BD9# else
		x"EE8A" when address_in = 16#0BDA# else
		x"EF9F" when address_in = 16#0BDB# else
		x"C013" when address_in = 16#0BDC# else
		x"835F" when address_in = 16#0BDD# else
		x"834E" when address_in = 16#0BDE# else
		x"838C" when address_in = 16#0BDF# else
		x"837B" when address_in = 16#0BE0# else
		x"836A" when address_in = 16#0BE1# else
		x"E082" when address_in = 16#0BE2# else
		x"838D" when address_in = 16#0BE3# else
		x"8219" when address_in = 16#0BE4# else
		x"8218" when address_in = 16#0BE5# else
		x"E020" when address_in = 16#0BE6# else
		x"E040" when address_in = 16#0BE7# else
		x"E050" when address_in = 16#0BE8# else
		x"2F8C" when address_in = 16#0BE9# else
		x"2F9D" when address_in = 16#0BEA# else
		x"940E" when address_in = 16#0BEB# else
		x"0B64" when address_in = 16#0BEC# else
		x"2799" when address_in = 16#0BED# else
		x"FD87" when address_in = 16#0BEE# else
		x"9590" when address_in = 16#0BEF# else
		x"91DF" when address_in = 16#0BF0# else
		x"91CF" when address_in = 16#0BF1# else
		x"9508" when address_in = 16#0BF2# else
		x"E786" when address_in = 16#0BF3# else
		x"E091" when address_in = 16#0BF4# else
		x"940E" when address_in = 16#0BF5# else
		x"116D" when address_in = 16#0BF6# else
		x"E083" when address_in = 16#0BF7# else
		x"E8E6" when address_in = 16#0BF8# else
		x"E0F1" when address_in = 16#0BF9# else
		x"9211" when address_in = 16#0BFA# else
		x"9211" when address_in = 16#0BFB# else
		x"5081" when address_in = 16#0BFC# else
		x"FF87" when address_in = 16#0BFD# else
		x"CFFB" when address_in = 16#0BFE# else
		x"EBE3" when address_in = 16#0BFF# else
		x"E0F0" when address_in = 16#0C00# else
		x"E083" when address_in = 16#0C01# else
		x"9211" when address_in = 16#0C02# else
		x"5081" when address_in = 16#0C03# else
		x"FF87" when address_in = 16#0C04# else
		x"CFFC" when address_in = 16#0C05# else
		x"E08E" when address_in = 16#0C06# else
		x"E099" when address_in = 16#0C07# else
		x"27AA" when address_in = 16#0C08# else
		x"FD97" when address_in = 16#0C09# else
		x"95A0" when address_in = 16#0C0A# else
		x"2FBA" when address_in = 16#0C0B# else
		x"95B6" when address_in = 16#0C0C# else
		x"95A7" when address_in = 16#0C0D# else
		x"9597" when address_in = 16#0C0E# else
		x"9587" when address_in = 16#0C0F# else
		x"E846" when address_in = 16#0C10# else
		x"E051" when address_in = 16#0C11# else
		x"2F68" when address_in = 16#0C12# else
		x"2F79" when address_in = 16#0C13# else
		x"E881" when address_in = 16#0C14# else
		x"E090" when address_in = 16#0C15# else
		x"940E" when address_in = 16#0C16# else
		x"0BC4" when address_in = 16#0C17# else
		x"E083" when address_in = 16#0C18# else
		x"E9E9" when address_in = 16#0C19# else
		x"E0F0" when address_in = 16#0C1A# else
		x"9211" when address_in = 16#0C1B# else
		x"9211" when address_in = 16#0C1C# else
		x"5081" when address_in = 16#0C1D# else
		x"FF87" when address_in = 16#0C1E# else
		x"CFFB" when address_in = 16#0C1F# else
		x"E889" when address_in = 16#0C20# else
		x"E090" when address_in = 16#0C21# else
		x"9390" when address_in = 16#0C22# else
		x"0175" when address_in = 16#0C23# else
		x"9380" when address_in = 16#0C24# else
		x"0174" when address_in = 16#0C25# else
		x"EA8D" when address_in = 16#0C26# else
		x"E090" when address_in = 16#0C27# else
		x"9390" when address_in = 16#0C28# else
		x"00AA" when address_in = 16#0C29# else
		x"9380" when address_in = 16#0C2A# else
		x"00A9" when address_in = 16#0C2B# else
		x"9180" when address_in = 16#0C2C# else
		x"0062" when address_in = 16#0C2D# else
		x"9190" when address_in = 16#0C2E# else
		x"0063" when address_in = 16#0C2F# else
		x"9390" when address_in = 16#0C30# else
		x"00A4" when address_in = 16#0C31# else
		x"9380" when address_in = 16#0C32# else
		x"00A3" when address_in = 16#0C33# else
		x"9390" when address_in = 16#0C34# else
		x"00A6" when address_in = 16#0C35# else
		x"9380" when address_in = 16#0C36# else
		x"00A5" when address_in = 16#0C37# else
		x"E083" when address_in = 16#0C38# else
		x"9380" when address_in = 16#0C39# else
		x"00A8" when address_in = 16#0C3A# else
		x"9508" when address_in = 16#0C3B# else
		x"92CF" when address_in = 16#0C3C# else
		x"92DF" when address_in = 16#0C3D# else
		x"92EF" when address_in = 16#0C3E# else
		x"92FF" when address_in = 16#0C3F# else
		x"930F" when address_in = 16#0C40# else
		x"931F" when address_in = 16#0C41# else
		x"93CF" when address_in = 16#0C42# else
		x"93DF" when address_in = 16#0C43# else
		x"2EE8" when address_in = 16#0C44# else
		x"2EF9" when address_in = 16#0C45# else
		x"2FD7" when address_in = 16#0C46# else
		x"2FC6" when address_in = 16#0C47# else
		x"2EC4" when address_in = 16#0C48# else
		x"2ED5" when address_in = 16#0C49# else
		x"2F12" when address_in = 16#0C4A# else
		x"3001" when address_in = 16#0C4B# else
		x"F521" when address_in = 16#0C4C# else
		x"E020" when address_in = 16#0C4D# else
		x"2F72" when address_in = 16#0C4E# else
		x"E031" when address_in = 16#0C4F# else
		x"E060" when address_in = 16#0C50# else
		x"2F47" when address_in = 16#0C51# else
		x"2755" when address_in = 16#0C52# else
		x"312F" when address_in = 16#0C53# else
		x"F081" when address_in = 16#0C54# else
		x"2FF5" when address_in = 16#0C55# else
		x"2FE4" when address_in = 16#0C56# else
		x"54ED" when address_in = 16#0C57# else
		x"4FFF" when address_in = 16#0C58# else
		x"8190" when address_in = 16#0C59# else
		x"2F83" when address_in = 16#0C5A# else
		x"2389" when address_in = 16#0C5B# else
		x"F071" when address_in = 16#0C5C# else
		x"5F6F" when address_in = 16#0C5D# else
		x"5F2F" when address_in = 16#0C5E# else
		x"0F33" when address_in = 16#0C5F# else
		x"3068" when address_in = 16#0C60# else
		x"F388" when address_in = 16#0C61# else
		x"5F7F" when address_in = 16#0C62# else
		x"3074" when address_in = 16#0C63# else
		x"F350" when address_in = 16#0C64# else
		x"EF8F" when address_in = 16#0C65# else
		x"E090" when address_in = 16#0C66# else
		x"2F08" when address_in = 16#0C67# else
		x"3F8F" when address_in = 16#0C68# else
		x"F4C9" when address_in = 16#0C69# else
		x"C032" when address_in = 16#0C6A# else
		x"2B93" when address_in = 16#0C6B# else
		x"8390" when address_in = 16#0C6C# else
		x"5220" when address_in = 16#0C6D# else
		x"2F82" when address_in = 16#0C6E# else
		x"2799" when address_in = 16#0C6F# else
		x"CFF6" when address_in = 16#0C70# else
		x"2D8E" when address_in = 16#0C71# else
		x"2D9F" when address_in = 16#0C72# else
		x"27AA" when address_in = 16#0C73# else
		x"27BB" when address_in = 16#0C74# else
		x"0F88" when address_in = 16#0C75# else
		x"1F99" when address_in = 16#0C76# else
		x"1FAA" when address_in = 16#0C77# else
		x"1FBB" when address_in = 16#0C78# else
		x"BFAB" when address_in = 16#0C79# else
		x"2FF9" when address_in = 16#0C7A# else
		x"2FE8" when address_in = 16#0C7B# else
		x"95D8" when address_in = 16#0C7C# else
		x"2D00" when address_in = 16#0C7D# else
		x"3E00" when address_in = 16#0C7E# else
		x"F018" when address_in = 16#0C7F# else
		x"EE8A" when address_in = 16#0C80# else
		x"EF9F" when address_in = 16#0C81# else
		x"C045" when address_in = 16#0C82# else
		x"2D8E" when address_in = 16#0C83# else
		x"2D9F" when address_in = 16#0C84# else
		x"27AA" when address_in = 16#0C85# else
		x"27BB" when address_in = 16#0C86# else
		x"0F88" when address_in = 16#0C87# else
		x"1F99" when address_in = 16#0C88# else
		x"1FAA" when address_in = 16#0C89# else
		x"1FBB" when address_in = 16#0C8A# else
		x"9601" when address_in = 16#0C8B# else
		x"1DA1" when address_in = 16#0C8C# else
		x"1DB1" when address_in = 16#0C8D# else
		x"BFAB" when address_in = 16#0C8E# else
		x"2FF9" when address_in = 16#0C8F# else
		x"2FE8" when address_in = 16#0C90# else
		x"95D8" when address_in = 16#0C91# else
		x"2D80" when address_in = 16#0C92# else
		x"2388" when address_in = 16#0C93# else
		x"F059" when address_in = 16#0C94# else
		x"E062" when address_in = 16#0C95# else
		x"2799" when address_in = 16#0C96# else
		x"940E" when address_in = 16#0C97# else
		x"0640" when address_in = 16#0C98# else
		x"839F" when address_in = 16#0C99# else
		x"838E" when address_in = 16#0C9A# else
		x"2B89" when address_in = 16#0C9B# else
		x"F429" when address_in = 16#0C9C# else
		x"EF84" when address_in = 16#0C9D# else
		x"EF9F" when address_in = 16#0C9E# else
		x"C028" when address_in = 16#0C9F# else
		x"821F" when address_in = 16#0CA0# else
		x"821E" when address_in = 16#0CA1# else
		x"82FB" when address_in = 16#0CA2# else
		x"82EA" when address_in = 16#0CA3# else
		x"830C" when address_in = 16#0CA4# else
		x"821D" when address_in = 16#0CA5# else
		x"8219" when address_in = 16#0CA6# else
		x"8218" when address_in = 16#0CA7# else
		x"2F21" when address_in = 16#0CA8# else
		x"2D5D" when address_in = 16#0CA9# else
		x"2D4C" when address_in = 16#0CAA# else
		x"2D7F" when address_in = 16#0CAB# else
		x"2D6E" when address_in = 16#0CAC# else
		x"2F8C" when address_in = 16#0CAD# else
		x"2F9D" when address_in = 16#0CAE# else
		x"940E" when address_in = 16#0CAF# else
		x"0B64" when address_in = 16#0CB0# else
		x"2F08" when address_in = 16#0CB1# else
		x"2388" when address_in = 16#0CB2# else
		x"F091" when address_in = 16#0CB3# else
		x"B184" when address_in = 16#0CB4# else
		x"2799" when address_in = 16#0CB5# else
		x"718E" when address_in = 16#0CB6# else
		x"7090" when address_in = 16#0CB7# else
		x"9595" when address_in = 16#0CB8# else
		x"9587" when address_in = 16#0CB9# else
		x"9595" when address_in = 16#0CBA# else
		x"9587" when address_in = 16#0CBB# else
		x"2F68" when address_in = 16#0CBC# else
		x"818E" when address_in = 16#0CBD# else
		x"819F" when address_in = 16#0CBE# else
		x"940E" when address_in = 16#0CBF# else
		x"07EC" when address_in = 16#0CC0# else
		x"2F80" when address_in = 16#0CC1# else
		x"2799" when address_in = 16#0CC2# else
		x"FD87" when address_in = 16#0CC3# else
		x"9590" when address_in = 16#0CC4# else
		x"C002" when address_in = 16#0CC5# else
		x"E080" when address_in = 16#0CC6# else
		x"E090" when address_in = 16#0CC7# else
		x"91DF" when address_in = 16#0CC8# else
		x"91CF" when address_in = 16#0CC9# else
		x"911F" when address_in = 16#0CCA# else
		x"910F" when address_in = 16#0CCB# else
		x"90FF" when address_in = 16#0CCC# else
		x"90EF" when address_in = 16#0CCD# else
		x"90DF" when address_in = 16#0CCE# else
		x"90CF" when address_in = 16#0CCF# else
		x"9508" when address_in = 16#0CD0# else
		x"92CF" when address_in = 16#0CD1# else
		x"92DF" when address_in = 16#0CD2# else
		x"92EF" when address_in = 16#0CD3# else
		x"92FF" when address_in = 16#0CD4# else
		x"930F" when address_in = 16#0CD5# else
		x"931F" when address_in = 16#0CD6# else
		x"93CF" when address_in = 16#0CD7# else
		x"93DF" when address_in = 16#0CD8# else
		x"2EE8" when address_in = 16#0CD9# else
		x"2EF9" when address_in = 16#0CDA# else
		x"2EC6" when address_in = 16#0CDB# else
		x"2ED7" when address_in = 16#0CDC# else
		x"2F14" when address_in = 16#0CDD# else
		x"2F02" when address_in = 16#0CDE# else
		x"2B89" when address_in = 16#0CDF# else
		x"F109" when address_in = 16#0CE0# else
		x"E062" when address_in = 16#0CE1# else
		x"E088" when address_in = 16#0CE2# else
		x"E090" when address_in = 16#0CE3# else
		x"940E" when address_in = 16#0CE4# else
		x"0640" when address_in = 16#0CE5# else
		x"2FD9" when address_in = 16#0CE6# else
		x"2FC8" when address_in = 16#0CE7# else
		x"9700" when address_in = 16#0CE8# else
		x"F0C1" when address_in = 16#0CE9# else
		x"2F21" when address_in = 16#0CEA# else
		x"2D5D" when address_in = 16#0CEB# else
		x"2D4C" when address_in = 16#0CEC# else
		x"2F68" when address_in = 16#0CED# else
		x"2F79" when address_in = 16#0CEE# else
		x"2D9F" when address_in = 16#0CEF# else
		x"2D8E" when address_in = 16#0CF0# else
		x"940E" when address_in = 16#0CF1# else
		x"0C3C" when address_in = 16#0CF2# else
		x"2388" when address_in = 16#0CF3# else
		x"F081" when address_in = 16#0CF4# else
		x"B184" when address_in = 16#0CF5# else
		x"2799" when address_in = 16#0CF6# else
		x"718E" when address_in = 16#0CF7# else
		x"7090" when address_in = 16#0CF8# else
		x"9595" when address_in = 16#0CF9# else
		x"9587" when address_in = 16#0CFA# else
		x"9595" when address_in = 16#0CFB# else
		x"9587" when address_in = 16#0CFC# else
		x"2F68" when address_in = 16#0CFD# else
		x"2F8C" when address_in = 16#0CFE# else
		x"2F9D" when address_in = 16#0CFF# else
		x"940E" when address_in = 16#0D00# else
		x"07EC" when address_in = 16#0D01# else
		x"EF8F" when address_in = 16#0D02# else
		x"E090" when address_in = 16#0D03# else
		x"C002" when address_in = 16#0D04# else
		x"818C" when address_in = 16#0D05# else
		x"2799" when address_in = 16#0D06# else
		x"91DF" when address_in = 16#0D07# else
		x"91CF" when address_in = 16#0D08# else
		x"911F" when address_in = 16#0D09# else
		x"910F" when address_in = 16#0D0A# else
		x"90FF" when address_in = 16#0D0B# else
		x"90EF" when address_in = 16#0D0C# else
		x"90DF" when address_in = 16#0D0D# else
		x"90CF" when address_in = 16#0D0E# else
		x"9508" when address_in = 16#0D0F# else
		x"92EF" when address_in = 16#0D10# else
		x"92FF" when address_in = 16#0D11# else
		x"930F" when address_in = 16#0D12# else
		x"93CF" when address_in = 16#0D13# else
		x"93DF" when address_in = 16#0D14# else
		x"2EE8" when address_in = 16#0D15# else
		x"2EF9" when address_in = 16#0D16# else
		x"2B89" when address_in = 16#0D17# else
		x"F419" when address_in = 16#0D18# else
		x"EE8A" when address_in = 16#0D19# else
		x"EF9F" when address_in = 16#0D1A# else
		x"C039" when address_in = 16#0D1B# else
		x"E062" when address_in = 16#0D1C# else
		x"E088" when address_in = 16#0D1D# else
		x"E090" when address_in = 16#0D1E# else
		x"940E" when address_in = 16#0D1F# else
		x"0640" when address_in = 16#0D20# else
		x"2FD9" when address_in = 16#0D21# else
		x"2FC8" when address_in = 16#0D22# else
		x"9700" when address_in = 16#0D23# else
		x"F419" when address_in = 16#0D24# else
		x"EF84" when address_in = 16#0D25# else
		x"EF9F" when address_in = 16#0D26# else
		x"C02D" when address_in = 16#0D27# else
		x"E000" when address_in = 16#0D28# else
		x"2F20" when address_in = 16#0D29# else
		x"E040" when address_in = 16#0D2A# else
		x"E050" when address_in = 16#0D2B# else
		x"2F68" when address_in = 16#0D2C# else
		x"2F79" when address_in = 16#0D2D# else
		x"2D9F" when address_in = 16#0D2E# else
		x"2D8E" when address_in = 16#0D2F# else
		x"940E" when address_in = 16#0D30# else
		x"0C3C" when address_in = 16#0D31# else
		x"2F08" when address_in = 16#0D32# else
		x"2388" when address_in = 16#0D33# else
		x"F069" when address_in = 16#0D34# else
		x"B184" when address_in = 16#0D35# else
		x"2799" when address_in = 16#0D36# else
		x"718E" when address_in = 16#0D37# else
		x"7090" when address_in = 16#0D38# else
		x"9595" when address_in = 16#0D39# else
		x"9587" when address_in = 16#0D3A# else
		x"9595" when address_in = 16#0D3B# else
		x"9587" when address_in = 16#0D3C# else
		x"2F68" when address_in = 16#0D3D# else
		x"2F8C" when address_in = 16#0D3E# else
		x"2F9D" when address_in = 16#0D3F# else
		x"940E" when address_in = 16#0D40# else
		x"07EC" when address_in = 16#0D41# else
		x"812C" when address_in = 16#0D42# else
		x"B184" when address_in = 16#0D43# else
		x"2799" when address_in = 16#0D44# else
		x"718E" when address_in = 16#0D45# else
		x"7090" when address_in = 16#0D46# else
		x"9595" when address_in = 16#0D47# else
		x"9587" when address_in = 16#0D48# else
		x"9595" when address_in = 16#0D49# else
		x"9587" when address_in = 16#0D4A# else
		x"2F48" when address_in = 16#0D4B# else
		x"2F62" when address_in = 16#0D4C# else
		x"818E" when address_in = 16#0D4D# else
		x"819F" when address_in = 16#0D4E# else
		x"940E" when address_in = 16#0D4F# else
		x"0700" when address_in = 16#0D50# else
		x"2F80" when address_in = 16#0D51# else
		x"2799" when address_in = 16#0D52# else
		x"FD87" when address_in = 16#0D53# else
		x"9590" when address_in = 16#0D54# else
		x"91DF" when address_in = 16#0D55# else
		x"91CF" when address_in = 16#0D56# else
		x"910F" when address_in = 16#0D57# else
		x"90FF" when address_in = 16#0D58# else
		x"90EF" when address_in = 16#0D59# else
		x"9508" when address_in = 16#0D5A# else
		x"92AF" when address_in = 16#0D5B# else
		x"92BF" when address_in = 16#0D5C# else
		x"92CF" when address_in = 16#0D5D# else
		x"92DF" when address_in = 16#0D5E# else
		x"92EF" when address_in = 16#0D5F# else
		x"92FF" when address_in = 16#0D60# else
		x"930F" when address_in = 16#0D61# else
		x"931F" when address_in = 16#0D62# else
		x"93CF" when address_in = 16#0D63# else
		x"93DF" when address_in = 16#0D64# else
		x"B7CD" when address_in = 16#0D65# else
		x"B7DE" when address_in = 16#0D66# else
		x"9762" when address_in = 16#0D67# else
		x"B60F" when address_in = 16#0D68# else
		x"94F8" when address_in = 16#0D69# else
		x"BFDE" when address_in = 16#0D6A# else
		x"BE0F" when address_in = 16#0D6B# else
		x"BFCD" when address_in = 16#0D6C# else
		x"2F08" when address_in = 16#0D6D# else
		x"7083" when address_in = 16#0D6E# else
		x"24AA" when address_in = 16#0D6F# else
		x"24BB" when address_in = 16#0D70# else
		x"2EC8" when address_in = 16#0D71# else
		x"24DD" when address_in = 16#0D72# else
		x"2DFD" when address_in = 16#0D73# else
		x"2DEC" when address_in = 16#0D74# else
		x"0DEC" when address_in = 16#0D75# else
		x"1DFD" when address_in = 16#0D76# else
		x"57EA" when address_in = 16#0D77# else
		x"4FFE" when address_in = 16#0D78# else
		x"80E0" when address_in = 16#0D79# else
		x"80F1" when address_in = 16#0D7A# else
		x"14E1" when address_in = 16#0D7B# else
		x"04F1" when address_in = 16#0D7C# else
		x"F041" when address_in = 16#0D7D# else
		x"2DFF" when address_in = 16#0D7E# else
		x"2DEE" when address_in = 16#0D7F# else
		x"8184" when address_in = 16#0D80# else
		x"1780" when address_in = 16#0D81# else
		x"F019" when address_in = 16#0D82# else
		x"2CAE" when address_in = 16#0D83# else
		x"2CBF" when address_in = 16#0D84# else
		x"CFF3" when address_in = 16#0D85# else
		x"14E1" when address_in = 16#0D86# else
		x"04F1" when address_in = 16#0D87# else
		x"F419" when address_in = 16#0D88# else
		x"EE8A" when address_in = 16#0D89# else
		x"EF9F" when address_in = 16#0D8A# else
		x"C08A" when address_in = 16#0D8B# else
		x"2DFF" when address_in = 16#0D8C# else
		x"2DEE" when address_in = 16#0D8D# else
		x"8182" when address_in = 16#0D8E# else
		x"8193" when address_in = 16#0D8F# else
		x"27AA" when address_in = 16#0D90# else
		x"27BB" when address_in = 16#0D91# else
		x"0F88" when address_in = 16#0D92# else
		x"1F99" when address_in = 16#0D93# else
		x"1FAA" when address_in = 16#0D94# else
		x"1FBB" when address_in = 16#0D95# else
		x"960C" when address_in = 16#0D96# else
		x"1DA1" when address_in = 16#0D97# else
		x"1DB1" when address_in = 16#0D98# else
		x"BFAB" when address_in = 16#0D99# else
		x"2FF9" when address_in = 16#0D9A# else
		x"2FE8" when address_in = 16#0D9B# else
		x"95D8" when address_in = 16#0D9C# else
		x"2D40" when address_in = 16#0D9D# else
		x"B60B" when address_in = 16#0D9E# else
		x"9631" when address_in = 16#0D9F# else
		x"1C01" when address_in = 16#0DA0# else
		x"BE0B" when address_in = 16#0DA1# else
		x"95D8" when address_in = 16#0DA2# else
		x"2D50" when address_in = 16#0DA3# else
		x"1541" when address_in = 16#0DA4# else
		x"0551" when address_in = 16#0DA5# else
		x"F0F9" when address_in = 16#0DA6# else
		x"2DFF" when address_in = 16#0DA7# else
		x"2DEE" when address_in = 16#0DA8# else
		x"8126" when address_in = 16#0DA9# else
		x"8137" when address_in = 16#0DAA# else
		x"9110" when address_in = 16#0DAB# else
		x"0173" when address_in = 16#0DAC# else
		x"8184" when address_in = 16#0DAD# else
		x"9380" when address_in = 16#0DAE# else
		x"0173" when address_in = 16#0DAF# else
		x"8184" when address_in = 16#0DB0# else
		x"8389" when address_in = 16#0DB1# else
		x"E082" when address_in = 16#0DB2# else
		x"838A" when address_in = 16#0DB3# else
		x"E086" when address_in = 16#0DB4# else
		x"838F" when address_in = 16#0DB5# else
		x"8618" when address_in = 16#0DB6# else
		x"861A" when address_in = 16#0DB7# else
		x"8619" when address_in = 16#0DB8# else
		x"861C" when address_in = 16#0DB9# else
		x"861B" when address_in = 16#0DBA# else
		x"2F6C" when address_in = 16#0DBB# else
		x"2F7D" when address_in = 16#0DBC# else
		x"5F6F" when address_in = 16#0DBD# else
		x"4F7F" when address_in = 16#0DBE# else
		x"2F93" when address_in = 16#0DBF# else
		x"2F82" when address_in = 16#0DC0# else
		x"2FE4" when address_in = 16#0DC1# else
		x"2FF5" when address_in = 16#0DC2# else
		x"9509" when address_in = 16#0DC3# else
		x"9310" when address_in = 16#0DC4# else
		x"0173" when address_in = 16#0DC5# else
		x"B72F" when address_in = 16#0DC6# else
		x"94F8" when address_in = 16#0DC7# else
		x"2DFF" when address_in = 16#0DC8# else
		x"2DEE" when address_in = 16#0DC9# else
		x"8180" when address_in = 16#0DCA# else
		x"8191" when address_in = 16#0DCB# else
		x"14A1" when address_in = 16#0DCC# else
		x"04B1" when address_in = 16#0DCD# else
		x"F449" when address_in = 16#0DCE# else
		x"0CCC" when address_in = 16#0DCF# else
		x"1CDD" when address_in = 16#0DD0# else
		x"E846" when address_in = 16#0DD1# else
		x"E051" when address_in = 16#0DD2# else
		x"0EC4" when address_in = 16#0DD3# else
		x"1ED5" when address_in = 16#0DD4# else
		x"2DFD" when address_in = 16#0DD5# else
		x"2DEC" when address_in = 16#0DD6# else
		x"C002" when address_in = 16#0DD7# else
		x"2DFB" when address_in = 16#0DD8# else
		x"2DEA" when address_in = 16#0DD9# else
		x"8391" when address_in = 16#0DDA# else
		x"8380" when address_in = 16#0DDB# else
		x"BF2F" when address_in = 16#0DDC# else
		x"2DFF" when address_in = 16#0DDD# else
		x"2DEE" when address_in = 16#0DDE# else
		x"8124" when address_in = 16#0DDF# else
		x"3E20" when address_in = 16#0DE0# else
		x"F0B0" when address_in = 16#0DE1# else
		x"5E20" when address_in = 16#0DE2# else
		x"2F82" when address_in = 16#0DE3# else
		x"9586" when address_in = 16#0DE4# else
		x"9586" when address_in = 16#0DE5# else
		x"9586" when address_in = 16#0DE6# else
		x"2FE8" when address_in = 16#0DE7# else
		x"27FF" when address_in = 16#0DE8# else
		x"54ED" when address_in = 16#0DE9# else
		x"4FFF" when address_in = 16#0DEA# else
		x"7027" when address_in = 16#0DEB# else
		x"E081" when address_in = 16#0DEC# else
		x"E090" when address_in = 16#0DED# else
		x"C002" when address_in = 16#0DEE# else
		x"0F88" when address_in = 16#0DEF# else
		x"1F99" when address_in = 16#0DF0# else
		x"952A" when address_in = 16#0DF1# else
		x"F7E2" when address_in = 16#0DF2# else
		x"2F98" when address_in = 16#0DF3# else
		x"9590" when address_in = 16#0DF4# else
		x"8180" when address_in = 16#0DF5# else
		x"2389" when address_in = 16#0DF6# else
		x"8380" when address_in = 16#0DF7# else
		x"2F80" when address_in = 16#0DF8# else
		x"940E" when address_in = 16#0DF9# else
		x"1BAF" when address_in = 16#0DFA# else
		x"2D9F" when address_in = 16#0DFB# else
		x"2D8E" when address_in = 16#0DFC# else
		x"940E" when address_in = 16#0DFD# else
		x"1A43" when address_in = 16#0DFE# else
		x"2DFF" when address_in = 16#0DFF# else
		x"2DEE" when address_in = 16#0E00# else
		x"8185" when address_in = 16#0E01# else
		x"FD81" when address_in = 16#0E02# else
		x"C00D" when address_in = 16#0E03# else
		x"B184" when address_in = 16#0E04# else
		x"2799" when address_in = 16#0E05# else
		x"718E" when address_in = 16#0E06# else
		x"7090" when address_in = 16#0E07# else
		x"9595" when address_in = 16#0E08# else
		x"9587" when address_in = 16#0E09# else
		x"9595" when address_in = 16#0E0A# else
		x"9587" when address_in = 16#0E0B# else
		x"2F68" when address_in = 16#0E0C# else
		x"2D9F" when address_in = 16#0E0D# else
		x"2D8E" when address_in = 16#0E0E# else
		x"940E" when address_in = 16#0E0F# else
		x"07EC" when address_in = 16#0E10# else
		x"2F80" when address_in = 16#0E11# else
		x"940E" when address_in = 16#0E12# else
		x"0942" when address_in = 16#0E13# else
		x"E080" when address_in = 16#0E14# else
		x"E090" when address_in = 16#0E15# else
		x"9662" when address_in = 16#0E16# else
		x"B60F" when address_in = 16#0E17# else
		x"94F8" when address_in = 16#0E18# else
		x"BFDE" when address_in = 16#0E19# else
		x"BE0F" when address_in = 16#0E1A# else
		x"BFCD" when address_in = 16#0E1B# else
		x"91DF" when address_in = 16#0E1C# else
		x"91CF" when address_in = 16#0E1D# else
		x"911F" when address_in = 16#0E1E# else
		x"910F" when address_in = 16#0E1F# else
		x"90FF" when address_in = 16#0E20# else
		x"90EF" when address_in = 16#0E21# else
		x"90DF" when address_in = 16#0E22# else
		x"90CF" when address_in = 16#0E23# else
		x"90BF" when address_in = 16#0E24# else
		x"90AF" when address_in = 16#0E25# else
		x"9508" when address_in = 16#0E26# else
		x"930F" when address_in = 16#0E27# else
		x"931F" when address_in = 16#0E28# else
		x"93CF" when address_in = 16#0E29# else
		x"93DF" when address_in = 16#0E2A# else
		x"2F08" when address_in = 16#0E2B# else
		x"2F19" when address_in = 16#0E2C# else
		x"E030" when address_in = 16#0E2D# else
		x"2F23" when address_in = 16#0E2E# else
		x"E846" when address_in = 16#0E2F# else
		x"E051" when address_in = 16#0E30# else
		x"2FF5" when address_in = 16#0E31# else
		x"2FE4" when address_in = 16#0E32# else
		x"91C1" when address_in = 16#0E33# else
		x"91D1" when address_in = 16#0E34# else
		x"2F4E" when address_in = 16#0E35# else
		x"2F5F" when address_in = 16#0E36# else
		x"9720" when address_in = 16#0E37# else
		x"F109" when address_in = 16#0E38# else
		x"818A" when address_in = 16#0E39# else
		x"819B" when address_in = 16#0E3A# else
		x"27AA" when address_in = 16#0E3B# else
		x"27BB" when address_in = 16#0E3C# else
		x"0F88" when address_in = 16#0E3D# else
		x"1F99" when address_in = 16#0E3E# else
		x"1FAA" when address_in = 16#0E3F# else
		x"1FBB" when address_in = 16#0E40# else
		x"9608" when address_in = 16#0E41# else
		x"1DA1" when address_in = 16#0E42# else
		x"1DB1" when address_in = 16#0E43# else
		x"BFAB" when address_in = 16#0E44# else
		x"2FF9" when address_in = 16#0E45# else
		x"2FE8" when address_in = 16#0E46# else
		x"95D8" when address_in = 16#0E47# else
		x"2D80" when address_in = 16#0E48# else
		x"B60B" when address_in = 16#0E49# else
		x"9631" when address_in = 16#0E4A# else
		x"1C01" when address_in = 16#0E4B# else
		x"BE0B" when address_in = 16#0E4C# else
		x"95D8" when address_in = 16#0E4D# else
		x"2D90" when address_in = 16#0E4E# else
		x"1780" when address_in = 16#0E4F# else
		x"0791" when address_in = 16#0E50# else
		x"F421" when address_in = 16#0E51# else
		x"818C" when address_in = 16#0E52# else
		x"940E" when address_in = 16#0E53# else
		x"0D5B" when address_in = 16#0E54# else
		x"CFD7" when address_in = 16#0E55# else
		x"9009" when address_in = 16#0E56# else
		x"81D8" when address_in = 16#0E57# else
		x"2DC0" when address_in = 16#0E58# else
		x"CFDD" when address_in = 16#0E59# else
		x"3031" when address_in = 16#0E5A# else
		x"F019" when address_in = 16#0E5B# else
		x"5F2F" when address_in = 16#0E5C# else
		x"3024" when address_in = 16#0E5D# else
		x"F290" when address_in = 16#0E5E# else
		x"3031" when address_in = 16#0E5F# else
		x"F409" when address_in = 16#0E60# else
		x"CFCB" when address_in = 16#0E61# else
		x"91DF" when address_in = 16#0E62# else
		x"91CF" when address_in = 16#0E63# else
		x"911F" when address_in = 16#0E64# else
		x"910F" when address_in = 16#0E65# else
		x"9508" when address_in = 16#0E66# else
		x"92AF" when address_in = 16#0E67# else
		x"92BF" when address_in = 16#0E68# else
		x"92CF" when address_in = 16#0E69# else
		x"92DF" when address_in = 16#0E6A# else
		x"92EF" when address_in = 16#0E6B# else
		x"92FF" when address_in = 16#0E6C# else
		x"930F" when address_in = 16#0E6D# else
		x"931F" when address_in = 16#0E6E# else
		x"93CF" when address_in = 16#0E6F# else
		x"93DF" when address_in = 16#0E70# else
		x"2ED8" when address_in = 16#0E71# else
		x"2EC6" when address_in = 16#0E72# else
		x"2EB4" when address_in = 16#0E73# else
		x"2EA2" when address_in = 16#0E74# else
		x"940E" when address_in = 16#0E75# else
		x"0B28" when address_in = 16#0E76# else
		x"2FD9" when address_in = 16#0E77# else
		x"2FC8" when address_in = 16#0E78# else
		x"2B89" when address_in = 16#0E79# else
		x"F181" when address_in = 16#0E7A# else
		x"818A" when address_in = 16#0E7B# else
		x"819B" when address_in = 16#0E7C# else
		x"27AA" when address_in = 16#0E7D# else
		x"27BB" when address_in = 16#0E7E# else
		x"0F88" when address_in = 16#0E7F# else
		x"1F99" when address_in = 16#0E80# else
		x"1FAA" when address_in = 16#0E81# else
		x"1FBB" when address_in = 16#0E82# else
		x"960C" when address_in = 16#0E83# else
		x"1DA1" when address_in = 16#0E84# else
		x"1DB1" when address_in = 16#0E85# else
		x"BFAB" when address_in = 16#0E86# else
		x"2FF9" when address_in = 16#0E87# else
		x"2FE8" when address_in = 16#0E88# else
		x"95D8" when address_in = 16#0E89# else
		x"2D20" when address_in = 16#0E8A# else
		x"B60B" when address_in = 16#0E8B# else
		x"9631" when address_in = 16#0E8C# else
		x"1C01" when address_in = 16#0E8D# else
		x"BE0B" when address_in = 16#0E8E# else
		x"95D8" when address_in = 16#0E8F# else
		x"2D30" when address_in = 16#0E90# else
		x"818E" when address_in = 16#0E91# else
		x"819F" when address_in = 16#0E92# else
		x"91E0" when address_in = 16#0E93# else
		x"00A9" when address_in = 16#0E94# else
		x"91F0" when address_in = 16#0E95# else
		x"00AA" when address_in = 16#0E96# else
		x"92D0" when address_in = 16#0E97# else
		x"00A1" when address_in = 16#0E98# else
		x"92C0" when address_in = 16#0E99# else
		x"00A2" when address_in = 16#0E9A# else
		x"92B0" when address_in = 16#0E9B# else
		x"00A7" when address_in = 16#0E9C# else
		x"82A0" when address_in = 16#0E9D# else
		x"8312" when address_in = 16#0E9E# else
		x"8301" when address_in = 16#0E9F# else
		x"92F0" when address_in = 16#0EA0# else
		x"00AC" when address_in = 16#0EA1# else
		x"92E0" when address_in = 16#0EA2# else
		x"00AB" when address_in = 16#0EA3# else
		x"92D0" when address_in = 16#0EA4# else
		x"0173" when address_in = 16#0EA5# else
		x"EA61" when address_in = 16#0EA6# else
		x"E070" when address_in = 16#0EA7# else
		x"2FE2" when address_in = 16#0EA8# else
		x"2FF3" when address_in = 16#0EA9# else
		x"9509" when address_in = 16#0EAA# else
		x"91DF" when address_in = 16#0EAB# else
		x"91CF" when address_in = 16#0EAC# else
		x"911F" when address_in = 16#0EAD# else
		x"910F" when address_in = 16#0EAE# else
		x"90FF" when address_in = 16#0EAF# else
		x"90EF" when address_in = 16#0EB0# else
		x"90DF" when address_in = 16#0EB1# else
		x"90CF" when address_in = 16#0EB2# else
		x"90BF" when address_in = 16#0EB3# else
		x"90AF" when address_in = 16#0EB4# else
		x"9508" when address_in = 16#0EB5# else
		x"940E" when address_in = 16#0EB6# else
		x"0B28" when address_in = 16#0EB7# else
		x"2B89" when address_in = 16#0EB8# else
		x"F419" when address_in = 16#0EB9# else
		x"EE8A" when address_in = 16#0EBA# else
		x"EF9F" when address_in = 16#0EBB# else
		x"9508" when address_in = 16#0EBC# else
		x"E080" when address_in = 16#0EBD# else
		x"E090" when address_in = 16#0EBE# else
		x"9508" when address_in = 16#0EBF# else
		x"93CF" when address_in = 16#0EC0# else
		x"93DF" when address_in = 16#0EC1# else
		x"2FD9" when address_in = 16#0EC2# else
		x"2FC8" when address_in = 16#0EC3# else
		x"858A" when address_in = 16#0EC4# else
		x"859B" when address_in = 16#0EC5# else
		x"FF82" when address_in = 16#0EC6# else
		x"C00E" when address_in = 16#0EC7# else
		x"B184" when address_in = 16#0EC8# else
		x"2799" when address_in = 16#0EC9# else
		x"718E" when address_in = 16#0ECA# else
		x"7090" when address_in = 16#0ECB# else
		x"9595" when address_in = 16#0ECC# else
		x"9587" when address_in = 16#0ECD# else
		x"9595" when address_in = 16#0ECE# else
		x"9587" when address_in = 16#0ECF# else
		x"2F48" when address_in = 16#0ED0# else
		x"E062" when address_in = 16#0ED1# else
		x"8588" when address_in = 16#0ED2# else
		x"8599" when address_in = 16#0ED3# else
		x"940E" when address_in = 16#0ED4# else
		x"0700" when address_in = 16#0ED5# else
		x"2F6C" when address_in = 16#0ED6# else
		x"2F7D" when address_in = 16#0ED7# else
		x"E786" when address_in = 16#0ED8# else
		x"E091" when address_in = 16#0ED9# else
		x"940E" when address_in = 16#0EDA# else
		x"1180" when address_in = 16#0EDB# else
		x"91DF" when address_in = 16#0EDC# else
		x"91CF" when address_in = 16#0EDD# else
		x"9508" when address_in = 16#0EDE# else
		x"93CF" when address_in = 16#0EDF# else
		x"93DF" when address_in = 16#0EE0# else
		x"2FD9" when address_in = 16#0EE1# else
		x"2FC8" when address_in = 16#0EE2# else
		x"2F6C" when address_in = 16#0EE3# else
		x"2F7D" when address_in = 16#0EE4# else
		x"E786" when address_in = 16#0EE5# else
		x"E091" when address_in = 16#0EE6# else
		x"940E" when address_in = 16#0EE7# else
		x"129C" when address_in = 16#0EE8# else
		x"9700" when address_in = 16#0EE9# else
		x"F019" when address_in = 16#0EEA# else
		x"940E" when address_in = 16#0EEB# else
		x"134D" when address_in = 16#0EEC# else
		x"CFF5" when address_in = 16#0EED# else
		x"91DF" when address_in = 16#0EEE# else
		x"91CF" when address_in = 16#0EEF# else
		x"9508" when address_in = 16#0EF0# else
		x"93CF" when address_in = 16#0EF1# else
		x"2FC6" when address_in = 16#0EF2# else
		x"940E" when address_in = 16#0EF3# else
		x"0B28" when address_in = 16#0EF4# else
		x"2FF9" when address_in = 16#0EF5# else
		x"2FE8" when address_in = 16#0EF6# else
		x"2B89" when address_in = 16#0EF7# else
		x"F419" when address_in = 16#0EF8# else
		x"EE8A" when address_in = 16#0EF9# else
		x"EF9F" when address_in = 16#0EFA# else
		x"C007" when address_in = 16#0EFB# else
		x"8185" when address_in = 16#0EFC# else
		x"708F" when address_in = 16#0EFD# else
		x"7FC0" when address_in = 16#0EFE# else
		x"2B8C" when address_in = 16#0EFF# else
		x"8385" when address_in = 16#0F00# else
		x"E080" when address_in = 16#0F01# else
		x"E090" when address_in = 16#0F02# else
		x"91CF" when address_in = 16#0F03# else
		x"9508" when address_in = 16#0F04# else
		x"93CF" when address_in = 16#0F05# else
		x"93DF" when address_in = 16#0F06# else
		x"2FD7" when address_in = 16#0F07# else
		x"2FC6" when address_in = 16#0F08# else
		x"940E" when address_in = 16#0F09# else
		x"0B28" when address_in = 16#0F0A# else
		x"2FF9" when address_in = 16#0F0B# else
		x"2FE8" when address_in = 16#0F0C# else
		x"2B89" when address_in = 16#0F0D# else
		x"F419" when address_in = 16#0F0E# else
		x"EE8A" when address_in = 16#0F0F# else
		x"EF9F" when address_in = 16#0F10# else
		x"C005" when address_in = 16#0F11# else
		x"8185" when address_in = 16#0F12# else
		x"7F80" when address_in = 16#0F13# else
		x"8388" when address_in = 16#0F14# else
		x"E080" when address_in = 16#0F15# else
		x"E090" when address_in = 16#0F16# else
		x"91DF" when address_in = 16#0F17# else
		x"91CF" when address_in = 16#0F18# else
		x"9508" when address_in = 16#0F19# else
		x"928F" when address_in = 16#0F1A# else
		x"929F" when address_in = 16#0F1B# else
		x"92AF" when address_in = 16#0F1C# else
		x"92BF" when address_in = 16#0F1D# else
		x"92CF" when address_in = 16#0F1E# else
		x"92DF" when address_in = 16#0F1F# else
		x"92EF" when address_in = 16#0F20# else
		x"92FF" when address_in = 16#0F21# else
		x"930F" when address_in = 16#0F22# else
		x"931F" when address_in = 16#0F23# else
		x"93CF" when address_in = 16#0F24# else
		x"93DF" when address_in = 16#0F25# else
		x"9478" when address_in = 16#0F26# else
		x"94F8" when address_in = 16#0F27# else
		x"9180" when address_in = 16#0F28# else
		x"0080" when address_in = 16#0F29# else
		x"2388" when address_in = 16#0F2A# else
		x"F091" when address_in = 16#0F2B# else
		x"9478" when address_in = 16#0F2C# else
		x"9210" when address_in = 16#0F2D# else
		x"0080" when address_in = 16#0F2E# else
		x"E013" when address_in = 16#0F2F# else
		x"E9C9" when address_in = 16#0F30# else
		x"E0D0" when address_in = 16#0F31# else
		x"81E8" when address_in = 16#0F32# else
		x"81F9" when address_in = 16#0F33# else
		x"9730" when address_in = 16#0F34# else
		x"F019" when address_in = 16#0F35# else
		x"8219" when address_in = 16#0F36# else
		x"8218" when address_in = 16#0F37# else
		x"9509" when address_in = 16#0F38# else
		x"5011" when address_in = 16#0F39# else
		x"9622" when address_in = 16#0F3A# else
		x"FF17" when address_in = 16#0F3B# else
		x"CFF5" when address_in = 16#0F3C# else
		x"CFE9" when address_in = 16#0F3D# else
		x"9180" when address_in = 16#0F3E# else
		x"0176" when address_in = 16#0F3F# else
		x"2388" when address_in = 16#0F40# else
		x"F409" when address_in = 16#0F41# else
		x"C093" when address_in = 16#0F42# else
		x"9478" when address_in = 16#0F43# else
		x"24AA" when address_in = 16#0F44# else
		x"24BB" when address_in = 16#0F45# else
		x"EF7F" when address_in = 16#0F46# else
		x"2E97" when address_in = 16#0F47# else
		x"E062" when address_in = 16#0F48# else
		x"2E86" when address_in = 16#0F49# else
		x"E786" when address_in = 16#0F4A# else
		x"E091" when address_in = 16#0F4B# else
		x"940E" when address_in = 16#0F4C# else
		x"11CE" when address_in = 16#0F4D# else
		x"2FD9" when address_in = 16#0F4E# else
		x"2FC8" when address_in = 16#0F4F# else
		x"8188" when address_in = 16#0F50# else
		x"940E" when address_in = 16#0F51# else
		x"0B28" when address_in = 16#0F52# else
		x"2F08" when address_in = 16#0F53# else
		x"2F19" when address_in = 16#0F54# else
		x"818E" when address_in = 16#0F55# else
		x"3083" when address_in = 16#0F56# else
		x"F411" when address_in = 16#0F57# else
		x"84A8" when address_in = 16#0F58# else
		x"84B9" when address_in = 16#0F59# else
		x"858A" when address_in = 16#0F5A# else
		x"859B" when address_in = 16#0F5B# else
		x"FD83" when address_in = 16#0F5C# else
		x"8099" when address_in = 16#0F5D# else
		x"2F8C" when address_in = 16#0F5E# else
		x"2F9D" when address_in = 16#0F5F# else
		x"940E" when address_in = 16#0F60# else
		x"2310" when address_in = 16#0F61# else
		x"1501" when address_in = 16#0F62# else
		x"0511" when address_in = 16#0F63# else
		x"F409" when address_in = 16#0F64# else
		x"C052" when address_in = 16#0F65# else
		x"854A" when address_in = 16#0F66# else
		x"855B" when address_in = 16#0F67# else
		x"FF50" when address_in = 16#0F68# else
		x"C012" when address_in = 16#0F69# else
		x"2FF1" when address_in = 16#0F6A# else
		x"2FE0" when address_in = 16#0F6B# else
		x"8185" when address_in = 16#0F6C# else
		x"FD86" when address_in = 16#0F6D# else
		x"C00D" when address_in = 16#0F6E# else
		x"812A" when address_in = 16#0F6F# else
		x"813B" when address_in = 16#0F70# else
		x"9180" when address_in = 16#0F71# else
		x"0062" when address_in = 16#0F72# else
		x"9190" when address_in = 16#0F73# else
		x"0063" when address_in = 16#0F74# else
		x"1728" when address_in = 16#0F75# else
		x"0739" when address_in = 16#0F76# else
		x"F021" when address_in = 16#0F77# else
		x"5F2F" when address_in = 16#0F78# else
		x"4F3F" when address_in = 16#0F79# else
		x"F009" when address_in = 16#0F7A# else
		x"C03C" when address_in = 16#0F7B# else
		x"2FF1" when address_in = 16#0F7C# else
		x"2FE0" when address_in = 16#0F7D# else
		x"8182" when address_in = 16#0F7E# else
		x"8193" when address_in = 16#0F7F# else
		x"27AA" when address_in = 16#0F80# else
		x"27BB" when address_in = 16#0F81# else
		x"0F88" when address_in = 16#0F82# else
		x"1F99" when address_in = 16#0F83# else
		x"1FAA" when address_in = 16#0F84# else
		x"1FBB" when address_in = 16#0F85# else
		x"960C" when address_in = 16#0F86# else
		x"1DA1" when address_in = 16#0F87# else
		x"1DB1" when address_in = 16#0F88# else
		x"BFAB" when address_in = 16#0F89# else
		x"2FF9" when address_in = 16#0F8A# else
		x"2FE8" when address_in = 16#0F8B# else
		x"95D8" when address_in = 16#0F8C# else
		x"2CC0" when address_in = 16#0F8D# else
		x"B60B" when address_in = 16#0F8E# else
		x"9631" when address_in = 16#0F8F# else
		x"1C01" when address_in = 16#0F90# else
		x"BE0B" when address_in = 16#0F91# else
		x"95D8" when address_in = 16#0F92# else
		x"2CD0" when address_in = 16#0F93# else
		x"2FF1" when address_in = 16#0F94# else
		x"2FE0" when address_in = 16#0F95# else
		x"80E6" when address_in = 16#0F96# else
		x"80F7" when address_in = 16#0F97# else
		x"FF42" when address_in = 16#0F98# else
		x"C00F" when address_in = 16#0F99# else
		x"8128" when address_in = 16#0F9A# else
		x"B184" when address_in = 16#0F9B# else
		x"2799" when address_in = 16#0F9C# else
		x"718E" when address_in = 16#0F9D# else
		x"7090" when address_in = 16#0F9E# else
		x"9595" when address_in = 16#0F9F# else
		x"9587" when address_in = 16#0FA0# else
		x"9595" when address_in = 16#0FA1# else
		x"9587" when address_in = 16#0FA2# else
		x"2F48" when address_in = 16#0FA3# else
		x"2F62" when address_in = 16#0FA4# else
		x"8588" when address_in = 16#0FA5# else
		x"8599" when address_in = 16#0FA6# else
		x"940E" when address_in = 16#0FA7# else
		x"0700" when address_in = 16#0FA8# else
		x"2FF1" when address_in = 16#0FA9# else
		x"2FE0" when address_in = 16#0FAA# else
		x"8184" when address_in = 16#0FAB# else
		x"9380" when address_in = 16#0FAC# else
		x"0173" when address_in = 16#0FAD# else
		x"2F6C" when address_in = 16#0FAE# else
		x"2F7D" when address_in = 16#0FAF# else
		x"2D9F" when address_in = 16#0FB0# else
		x"2D8E" when address_in = 16#0FB1# else
		x"2DEC" when address_in = 16#0FB2# else
		x"2DFD" when address_in = 16#0FB3# else
		x"9509" when address_in = 16#0FB4# else
		x"2388" when address_in = 16#0FB5# else
		x"F409" when address_in = 16#0FB6# else
		x"2E88" when address_in = 16#0FB7# else
		x"14A1" when address_in = 16#0FB8# else
		x"04B1" when address_in = 16#0FB9# else
		x"F029" when address_in = 16#0FBA# else
		x"2D9B" when address_in = 16#0FBB# else
		x"2D8A" when address_in = 16#0FBC# else
		x"940E" when address_in = 16#0FBD# else
		x"134D" when address_in = 16#0FBE# else
		x"C011" when address_in = 16#0FBF# else
		x"EFFF" when address_in = 16#0FC0# else
		x"169F" when address_in = 16#0FC1# else
		x"F071" when address_in = 16#0FC2# else
		x"2D88" when address_in = 16#0FC3# else
		x"2799" when address_in = 16#0FC4# else
		x"2EE8" when address_in = 16#0FC5# else
		x"2EF9" when address_in = 16#0FC6# else
		x"2F0C" when address_in = 16#0FC7# else
		x"2F1D" when address_in = 16#0FC8# else
		x"E122" when address_in = 16#0FC9# else
		x"E043" when address_in = 16#0FCA# else
		x"E062" when address_in = 16#0FCB# else
		x"2D89" when address_in = 16#0FCC# else
		x"940E" when address_in = 16#0FCD# else
		x"105C" when address_in = 16#0FCE# else
		x"FF87" when address_in = 16#0FCF# else
		x"CF56" when address_in = 16#0FD0# else
		x"2F8C" when address_in = 16#0FD1# else
		x"2F9D" when address_in = 16#0FD2# else
		x"940E" when address_in = 16#0FD3# else
		x"134D" when address_in = 16#0FD4# else
		x"CF51" when address_in = 16#0FD5# else
		x"9478" when address_in = 16#0FD6# else
		x"CF4F" when address_in = 16#0FD7# else
		x"92BF" when address_in = 16#0FD8# else
		x"92CF" when address_in = 16#0FD9# else
		x"92DF" when address_in = 16#0FDA# else
		x"92EF" when address_in = 16#0FDB# else
		x"92FF" when address_in = 16#0FDC# else
		x"930F" when address_in = 16#0FDD# else
		x"931F" when address_in = 16#0FDE# else
		x"93CF" when address_in = 16#0FDF# else
		x"2ED8" when address_in = 16#0FE0# else
		x"2EC6" when address_in = 16#0FE1# else
		x"2FC4" when address_in = 16#0FE2# else
		x"2EB2" when address_in = 16#0FE3# else
		x"940E" when address_in = 16#0FE4# else
		x"12DE" when address_in = 16#0FE5# else
		x"2FF9" when address_in = 16#0FE6# else
		x"2FE8" when address_in = 16#0FE7# else
		x"2B89" when address_in = 16#0FE8# else
		x"F419" when address_in = 16#0FE9# else
		x"EF84" when address_in = 16#0FEA# else
		x"EF9F" when address_in = 16#0FEB# else
		x"C01F" when address_in = 16#0FEC# else
		x"9180" when address_in = 16#0FED# else
		x"0062" when address_in = 16#0FEE# else
		x"9190" when address_in = 16#0FEF# else
		x"0063" when address_in = 16#0FF0# else
		x"8393" when address_in = 16#0FF1# else
		x"8382" when address_in = 16#0FF2# else
		x"82D0" when address_in = 16#0FF3# else
		x"83C6" when address_in = 16#0FF4# else
		x"9180" when address_in = 16#0FF5# else
		x"0062" when address_in = 16#0FF6# else
		x"9190" when address_in = 16#0FF7# else
		x"0063" when address_in = 16#0FF8# else
		x"8395" when address_in = 16#0FF9# else
		x"8384" when address_in = 16#0FFA# else
		x"82C1" when address_in = 16#0FFB# else
		x"E083" when address_in = 16#0FFC# else
		x"8387" when address_in = 16#0FFD# else
		x"86B4" when address_in = 16#0FFE# else
		x"8716" when address_in = 16#0FFF# else
		x"8705" when address_in = 16#1000# else
		x"EF8B" when address_in = 16#1001# else
		x"22E8" when address_in = 16#1002# else
		x"24FF" when address_in = 16#1003# else
		x"86F3" when address_in = 16#1004# else
		x"86E2" when address_in = 16#1005# else
		x"2F8E" when address_in = 16#1006# else
		x"2F9F" when address_in = 16#1007# else
		x"940E" when address_in = 16#1008# else
		x"0EC0" when address_in = 16#1009# else
		x"E080" when address_in = 16#100A# else
		x"E090" when address_in = 16#100B# else
		x"91CF" when address_in = 16#100C# else
		x"911F" when address_in = 16#100D# else
		x"910F" when address_in = 16#100E# else
		x"90FF" when address_in = 16#100F# else
		x"90EF" when address_in = 16#1010# else
		x"90DF" when address_in = 16#1011# else
		x"90CF" when address_in = 16#1012# else
		x"90BF" when address_in = 16#1013# else
		x"9508" when address_in = 16#1014# else
		x"929F" when address_in = 16#1015# else
		x"92AF" when address_in = 16#1016# else
		x"92BF" when address_in = 16#1017# else
		x"92CF" when address_in = 16#1018# else
		x"92DF" when address_in = 16#1019# else
		x"92EF" when address_in = 16#101A# else
		x"92FF" when address_in = 16#101B# else
		x"930F" when address_in = 16#101C# else
		x"931F" when address_in = 16#101D# else
		x"93CF" when address_in = 16#101E# else
		x"2EB8" when address_in = 16#101F# else
		x"2E96" when address_in = 16#1020# else
		x"2FC4" when address_in = 16#1021# else
		x"2EA2" when address_in = 16#1022# else
		x"940E" when address_in = 16#1023# else
		x"12DE" when address_in = 16#1024# else
		x"2FF9" when address_in = 16#1025# else
		x"2FE8" when address_in = 16#1026# else
		x"2B89" when address_in = 16#1027# else
		x"F491" when address_in = 16#1028# else
		x"FEE2" when address_in = 16#1029# else
		x"C00D" when address_in = 16#102A# else
		x"B184" when address_in = 16#102B# else
		x"2799" when address_in = 16#102C# else
		x"718E" when address_in = 16#102D# else
		x"7090" when address_in = 16#102E# else
		x"9595" when address_in = 16#102F# else
		x"9587" when address_in = 16#1030# else
		x"9595" when address_in = 16#1031# else
		x"9587" when address_in = 16#1032# else
		x"2F68" when address_in = 16#1033# else
		x"2F91" when address_in = 16#1034# else
		x"2F80" when address_in = 16#1035# else
		x"940E" when address_in = 16#1036# else
		x"07EC" when address_in = 16#1037# else
		x"EF84" when address_in = 16#1038# else
		x"EF9F" when address_in = 16#1039# else
		x"C016" when address_in = 16#103A# else
		x"9180" when address_in = 16#103B# else
		x"0062" when address_in = 16#103C# else
		x"9190" when address_in = 16#103D# else
		x"0063" when address_in = 16#103E# else
		x"8393" when address_in = 16#103F# else
		x"8382" when address_in = 16#1040# else
		x"82B0" when address_in = 16#1041# else
		x"83C6" when address_in = 16#1042# else
		x"82D5" when address_in = 16#1043# else
		x"82C4" when address_in = 16#1044# else
		x"8291" when address_in = 16#1045# else
		x"82A7" when address_in = 16#1046# else
		x"8711" when address_in = 16#1047# else
		x"8700" when address_in = 16#1048# else
		x"86F3" when address_in = 16#1049# else
		x"86E2" when address_in = 16#104A# else
		x"2F8E" when address_in = 16#104B# else
		x"2F9F" when address_in = 16#104C# else
		x"940E" when address_in = 16#104D# else
		x"0EC0" when address_in = 16#104E# else
		x"E080" when address_in = 16#104F# else
		x"E090" when address_in = 16#1050# else
		x"91CF" when address_in = 16#1051# else
		x"911F" when address_in = 16#1052# else
		x"910F" when address_in = 16#1053# else
		x"90FF" when address_in = 16#1054# else
		x"90EF" when address_in = 16#1055# else
		x"90DF" when address_in = 16#1056# else
		x"90CF" when address_in = 16#1057# else
		x"90BF" when address_in = 16#1058# else
		x"90AF" when address_in = 16#1059# else
		x"909F" when address_in = 16#105A# else
		x"9508" when address_in = 16#105B# else
		x"92CF" when address_in = 16#105C# else
		x"92DF" when address_in = 16#105D# else
		x"92EF" when address_in = 16#105E# else
		x"92FF" when address_in = 16#105F# else
		x"930F" when address_in = 16#1060# else
		x"931F" when address_in = 16#1061# else
		x"2F76" when address_in = 16#1062# else
		x"2F64" when address_in = 16#1063# else
		x"2F92" when address_in = 16#1064# else
		x"90C0" when address_in = 16#1065# else
		x"0062" when address_in = 16#1066# else
		x"90D0" when address_in = 16#1067# else
		x"0063" when address_in = 16#1068# else
		x"2F29" when address_in = 16#1069# else
		x"2F46" when address_in = 16#106A# else
		x"2F67" when address_in = 16#106B# else
		x"940E" when address_in = 16#106C# else
		x"1015" when address_in = 16#106D# else
		x"2799" when address_in = 16#106E# else
		x"FD87" when address_in = 16#106F# else
		x"9590" when address_in = 16#1070# else
		x"911F" when address_in = 16#1071# else
		x"910F" when address_in = 16#1072# else
		x"90FF" when address_in = 16#1073# else
		x"90EF" when address_in = 16#1074# else
		x"90DF" when address_in = 16#1075# else
		x"90CF" when address_in = 16#1076# else
		x"9508" when address_in = 16#1077# else
		x"929F" when address_in = 16#1078# else
		x"92AF" when address_in = 16#1079# else
		x"92BF" when address_in = 16#107A# else
		x"92CF" when address_in = 16#107B# else
		x"92DF" when address_in = 16#107C# else
		x"92EF" when address_in = 16#107D# else
		x"92FF" when address_in = 16#107E# else
		x"930F" when address_in = 16#107F# else
		x"931F" when address_in = 16#1080# else
		x"93CF" when address_in = 16#1081# else
		x"2E98" when address_in = 16#1082# else
		x"2EA6" when address_in = 16#1083# else
		x"2EB4" when address_in = 16#1084# else
		x"2EC2" when address_in = 16#1085# else
		x"2ED3" when address_in = 16#1086# else
		x"940E" when address_in = 16#1087# else
		x"0B5D" when address_in = 16#1088# else
		x"2FC8" when address_in = 16#1089# else
		x"2EE0" when address_in = 16#108A# else
		x"2EF1" when address_in = 16#108B# else
		x"2D1D" when address_in = 16#108C# else
		x"2D0C" when address_in = 16#108D# else
		x"2D2B" when address_in = 16#108E# else
		x"2D4A" when address_in = 16#108F# else
		x"2F68" when address_in = 16#1090# else
		x"2D89" when address_in = 16#1091# else
		x"940E" when address_in = 16#1092# else
		x"105C" when address_in = 16#1093# else
		x"2388" when address_in = 16#1094# else
		x"F039" when address_in = 16#1095# else
		x"2F8C" when address_in = 16#1096# else
		x"940E" when address_in = 16#1097# else
		x"09FA" when address_in = 16#1098# else
		x"2799" when address_in = 16#1099# else
		x"FD87" when address_in = 16#109A# else
		x"9590" when address_in = 16#109B# else
		x"C002" when address_in = 16#109C# else
		x"E080" when address_in = 16#109D# else
		x"E090" when address_in = 16#109E# else
		x"91CF" when address_in = 16#109F# else
		x"911F" when address_in = 16#10A0# else
		x"910F" when address_in = 16#10A1# else
		x"90FF" when address_in = 16#10A2# else
		x"90EF" when address_in = 16#10A3# else
		x"90DF" when address_in = 16#10A4# else
		x"90CF" when address_in = 16#10A5# else
		x"90BF" when address_in = 16#10A6# else
		x"90AF" when address_in = 16#10A7# else
		x"909F" when address_in = 16#10A8# else
		x"9508" when address_in = 16#10A9# else
		x"930F" when address_in = 16#10AA# else
		x"931F" when address_in = 16#10AB# else
		x"93CF" when address_in = 16#10AC# else
		x"93DF" when address_in = 16#10AD# else
		x"2F38" when address_in = 16#10AE# else
		x"2FF7" when address_in = 16#10AF# else
		x"2FE6" when address_in = 16#10B0# else
		x"8186" when address_in = 16#10B1# else
		x"3083" when address_in = 16#10B2# else
		x"F419" when address_in = 16#10B3# else
		x"85C0" when address_in = 16#10B4# else
		x"85D1" when address_in = 16#10B5# else
		x"C002" when address_in = 16#10B6# else
		x"2FD7" when address_in = 16#10B7# else
		x"2FC6" when address_in = 16#10B8# else
		x"858A" when address_in = 16#10B9# else
		x"859B" when address_in = 16#10BA# else
		x"FF82" when address_in = 16#10BB# else
		x"C019" when address_in = 16#10BC# else
		x"B184" when address_in = 16#10BD# else
		x"2799" when address_in = 16#10BE# else
		x"718E" when address_in = 16#10BF# else
		x"7090" when address_in = 16#10C0# else
		x"9595" when address_in = 16#10C1# else
		x"9587" when address_in = 16#10C2# else
		x"9595" when address_in = 16#10C3# else
		x"9587" when address_in = 16#10C4# else
		x"2F48" when address_in = 16#10C5# else
		x"2F63" when address_in = 16#10C6# else
		x"8588" when address_in = 16#10C7# else
		x"8599" when address_in = 16#10C8# else
		x"940E" when address_in = 16#10C9# else
		x"0700" when address_in = 16#10CA# else
		x"8508" when address_in = 16#10CB# else
		x"8519" when address_in = 16#10CC# else
		x"821F" when address_in = 16#10CD# else
		x"8619" when address_in = 16#10CE# else
		x"8618" when address_in = 16#10CF# else
		x"858A" when address_in = 16#10D0# else
		x"859B" when address_in = 16#10D1# else
		x"7F8B" when address_in = 16#10D2# else
		x"879B" when address_in = 16#10D3# else
		x"878A" when address_in = 16#10D4# else
		x"C01F" when address_in = 16#10D5# else
		x"812F" when address_in = 16#10D6# else
		x"B184" when address_in = 16#10D7# else
		x"2799" when address_in = 16#10D8# else
		x"718E" when address_in = 16#10D9# else
		x"7090" when address_in = 16#10DA# else
		x"9595" when address_in = 16#10DB# else
		x"9587" when address_in = 16#10DC# else
		x"9595" when address_in = 16#10DD# else
		x"9587" when address_in = 16#10DE# else
		x"2F48" when address_in = 16#10DF# else
		x"2F63" when address_in = 16#10E0# else
		x"2F82" when address_in = 16#10E1# else
		x"2799" when address_in = 16#10E2# else
		x"940E" when address_in = 16#10E3# else
		x"0889" when address_in = 16#10E4# else
		x"2F08" when address_in = 16#10E5# else
		x"2F19" when address_in = 16#10E6# else
		x"2B89" when address_in = 16#10E7# else
		x"F061" when address_in = 16#10E8# else
		x"818F" when address_in = 16#10E9# else
		x"2799" when address_in = 16#10EA# else
		x"8528" when address_in = 16#10EB# else
		x"8539" when address_in = 16#10EC# else
		x"2F48" when address_in = 16#10ED# else
		x"2F59" when address_in = 16#10EE# else
		x"2F73" when address_in = 16#10EF# else
		x"2F62" when address_in = 16#10F0# else
		x"2F91" when address_in = 16#10F1# else
		x"2F80" when address_in = 16#10F2# else
		x"940E" when address_in = 16#10F3# else
		x"2E67" when address_in = 16#10F4# else
		x"2F91" when address_in = 16#10F5# else
		x"2F80" when address_in = 16#10F6# else
		x"91DF" when address_in = 16#10F7# else
		x"91CF" when address_in = 16#10F8# else
		x"911F" when address_in = 16#10F9# else
		x"910F" when address_in = 16#10FA# else
		x"9508" when address_in = 16#10FB# else
		x"92FF" when address_in = 16#10FC# else
		x"930F" when address_in = 16#10FD# else
		x"931F" when address_in = 16#10FE# else
		x"93CF" when address_in = 16#10FF# else
		x"93DF" when address_in = 16#1100# else
		x"2F08" when address_in = 16#1101# else
		x"2F19" when address_in = 16#1102# else
		x"940E" when address_in = 16#1103# else
		x"0B5D" when address_in = 16#1104# else
		x"2EF8" when address_in = 16#1105# else
		x"2F71" when address_in = 16#1106# else
		x"2F60" when address_in = 16#1107# else
		x"940E" when address_in = 16#1108# else
		x"10AA" when address_in = 16#1109# else
		x"2FD9" when address_in = 16#110A# else
		x"2FC8" when address_in = 16#110B# else
		x"2B89" when address_in = 16#110C# else
		x"F419" when address_in = 16#110D# else
		x"2D8F" when address_in = 16#110E# else
		x"940E" when address_in = 16#110F# else
		x"09FA" when address_in = 16#1110# else
		x"2F8C" when address_in = 16#1111# else
		x"2F9D" when address_in = 16#1112# else
		x"91DF" when address_in = 16#1113# else
		x"91CF" when address_in = 16#1114# else
		x"911F" when address_in = 16#1115# else
		x"910F" when address_in = 16#1116# else
		x"90FF" when address_in = 16#1117# else
		x"9508" when address_in = 16#1118# else
		x"92AF" when address_in = 16#1119# else
		x"92BF" when address_in = 16#111A# else
		x"92CF" when address_in = 16#111B# else
		x"92DF" when address_in = 16#111C# else
		x"92EF" when address_in = 16#111D# else
		x"92FF" when address_in = 16#111E# else
		x"930F" when address_in = 16#111F# else
		x"931F" when address_in = 16#1120# else
		x"93CF" when address_in = 16#1121# else
		x"93DF" when address_in = 16#1122# else
		x"2EB8" when address_in = 16#1123# else
		x"2EA6" when address_in = 16#1124# else
		x"2EC2" when address_in = 16#1125# else
		x"2ED3" when address_in = 16#1126# else
		x"2EE4" when address_in = 16#1127# else
		x"2EF5" when address_in = 16#1128# else
		x"940E" when address_in = 16#1129# else
		x"12DE" when address_in = 16#112A# else
		x"2FD9" when address_in = 16#112B# else
		x"2FC8" when address_in = 16#112C# else
		x"940E" when address_in = 16#112D# else
		x"0B5D" when address_in = 16#112E# else
		x"2F28" when address_in = 16#112F# else
		x"9720" when address_in = 16#1130# else
		x"F431" when address_in = 16#1131# else
		x"940E" when address_in = 16#1132# else
		x"09FA" when address_in = 16#1133# else
		x"2799" when address_in = 16#1134# else
		x"FD87" when address_in = 16#1135# else
		x"9590" when address_in = 16#1136# else
		x"C021" when address_in = 16#1137# else
		x"9180" when address_in = 16#1138# else
		x"0062" when address_in = 16#1139# else
		x"9190" when address_in = 16#113A# else
		x"0063" when address_in = 16#113B# else
		x"839B" when address_in = 16#113C# else
		x"838A" when address_in = 16#113D# else
		x"82B8" when address_in = 16#113E# else
		x"82AE" when address_in = 16#113F# else
		x"9180" when address_in = 16#1140# else
		x"0062" when address_in = 16#1141# else
		x"9190" when address_in = 16#1142# else
		x"0063" when address_in = 16#1143# else
		x"839D" when address_in = 16#1144# else
		x"838C" when address_in = 16#1145# else
		x"8329" when address_in = 16#1146# else
		x"E084" when address_in = 16#1147# else
		x"838F" when address_in = 16#1148# else
		x"85E8" when address_in = 16#1149# else
		x"85F9" when address_in = 16#114A# else
		x"82C0" when address_in = 16#114B# else
		x"82D1" when address_in = 16#114C# else
		x"82E2" when address_in = 16#114D# else
		x"82F3" when address_in = 16#114E# else
		x"7F0B" when address_in = 16#114F# else
		x"7010" when address_in = 16#1150# else
		x"871B" when address_in = 16#1151# else
		x"870A" when address_in = 16#1152# else
		x"2F8C" when address_in = 16#1153# else
		x"2F9D" when address_in = 16#1154# else
		x"940E" when address_in = 16#1155# else
		x"0EC0" when address_in = 16#1156# else
		x"E080" when address_in = 16#1157# else
		x"E090" when address_in = 16#1158# else
		x"91DF" when address_in = 16#1159# else
		x"91CF" when address_in = 16#115A# else
		x"911F" when address_in = 16#115B# else
		x"910F" when address_in = 16#115C# else
		x"90FF" when address_in = 16#115D# else
		x"90EF" when address_in = 16#115E# else
		x"90DF" when address_in = 16#115F# else
		x"90CF" when address_in = 16#1160# else
		x"90BF" when address_in = 16#1161# else
		x"90AF" when address_in = 16#1162# else
		x"9508" when address_in = 16#1163# else
		x"9210" when address_in = 16#1164# else
		x"00B8" when address_in = 16#1165# else
		x"9210" when address_in = 16#1166# else
		x"00B7" when address_in = 16#1167# else
		x"9210" when address_in = 16#1168# else
		x"0101" when address_in = 16#1169# else
		x"E080" when address_in = 16#116A# else
		x"E090" when address_in = 16#116B# else
		x"9508" when address_in = 16#116C# else
		x"2FF9" when address_in = 16#116D# else
		x"2FE8" when address_in = 16#116E# else
		x"8210" when address_in = 16#116F# else
		x"8213" when address_in = 16#1170# else
		x"8212" when address_in = 16#1171# else
		x"8211" when address_in = 16#1172# else
		x"8215" when address_in = 16#1173# else
		x"8214" when address_in = 16#1174# else
		x"8217" when address_in = 16#1175# else
		x"8216" when address_in = 16#1176# else
		x"8611" when address_in = 16#1177# else
		x"8610" when address_in = 16#1178# else
		x"8613" when address_in = 16#1179# else
		x"8612" when address_in = 16#117A# else
		x"8615" when address_in = 16#117B# else
		x"8614" when address_in = 16#117C# else
		x"8617" when address_in = 16#117D# else
		x"8616" when address_in = 16#117E# else
		x"9508" when address_in = 16#117F# else
		x"93CF" when address_in = 16#1180# else
		x"93DF" when address_in = 16#1181# else
		x"2FD9" when address_in = 16#1182# else
		x"2FC8" when address_in = 16#1183# else
		x"2FB7" when address_in = 16#1184# else
		x"2FA6" when address_in = 16#1185# else
		x"B72F" when address_in = 16#1186# else
		x"94F8" when address_in = 16#1187# else
		x"2FF7" when address_in = 16#1188# else
		x"2FE6" when address_in = 16#1189# else
		x"8A11" when address_in = 16#118A# else
		x"8A10" when address_in = 16#118B# else
		x"8582" when address_in = 16#118C# else
		x"8593" when address_in = 16#118D# else
		x"FF86" when address_in = 16#118E# else
		x"C011" when address_in = 16#118F# else
		x"818C" when address_in = 16#1190# else
		x"819D" when address_in = 16#1191# else
		x"2B89" when address_in = 16#1192# else
		x"F419" when address_in = 16#1193# else
		x"837D" when address_in = 16#1194# else
		x"836C" when address_in = 16#1195# else
		x"C004" when address_in = 16#1196# else
		x"81EE" when address_in = 16#1197# else
		x"81FF" when address_in = 16#1198# else
		x"8B71" when address_in = 16#1199# else
		x"8B60" when address_in = 16#119A# else
		x"83BF" when address_in = 16#119B# else
		x"83AE" when address_in = 16#119C# else
		x"818B" when address_in = 16#119D# else
		x"5F8F" when address_in = 16#119E# else
		x"838B" when address_in = 16#119F# else
		x"C026" when address_in = 16#11A0# else
		x"2FF7" when address_in = 16#11A1# else
		x"2FE6" when address_in = 16#11A2# else
		x"8582" when address_in = 16#11A3# else
		x"FF87" when address_in = 16#11A4# else
		x"C011" when address_in = 16#11A5# else
		x"8588" when address_in = 16#11A6# else
		x"8599" when address_in = 16#11A7# else
		x"2B89" when address_in = 16#11A8# else
		x"F419" when address_in = 16#11A9# else
		x"8779" when address_in = 16#11AA# else
		x"8768" when address_in = 16#11AB# else
		x"C004" when address_in = 16#11AC# else
		x"85EA" when address_in = 16#11AD# else
		x"85FB" when address_in = 16#11AE# else
		x"8B71" when address_in = 16#11AF# else
		x"8B60" when address_in = 16#11B0# else
		x"87BB" when address_in = 16#11B1# else
		x"87AA" when address_in = 16#11B2# else
		x"818A" when address_in = 16#11B3# else
		x"5F8F" when address_in = 16#11B4# else
		x"838A" when address_in = 16#11B5# else
		x"C010" when address_in = 16#11B6# else
		x"858C" when address_in = 16#11B7# else
		x"859D" when address_in = 16#11B8# else
		x"2B89" when address_in = 16#11B9# else
		x"F419" when address_in = 16#11BA# else
		x"877D" when address_in = 16#11BB# else
		x"876C" when address_in = 16#11BC# else
		x"C004" when address_in = 16#11BD# else
		x"85EE" when address_in = 16#11BE# else
		x"85FF" when address_in = 16#11BF# else
		x"8B71" when address_in = 16#11C0# else
		x"8B60" when address_in = 16#11C1# else
		x"87BF" when address_in = 16#11C2# else
		x"87AE" when address_in = 16#11C3# else
		x"8189" when address_in = 16#11C4# else
		x"5F8F" when address_in = 16#11C5# else
		x"8389" when address_in = 16#11C6# else
		x"8188" when address_in = 16#11C7# else
		x"5F8F" when address_in = 16#11C8# else
		x"8388" when address_in = 16#11C9# else
		x"BF2F" when address_in = 16#11CA# else
		x"91DF" when address_in = 16#11CB# else
		x"91CF" when address_in = 16#11CC# else
		x"9508" when address_in = 16#11CD# else
		x"93CF" when address_in = 16#11CE# else
		x"93DF" when address_in = 16#11CF# else
		x"2FF9" when address_in = 16#11D0# else
		x"2FE8" when address_in = 16#11D1# else
		x"B72F" when address_in = 16#11D2# else
		x"94F8" when address_in = 16#11D3# else
		x"81A4" when address_in = 16#11D4# else
		x"81B5" when address_in = 16#11D5# else
		x"9710" when address_in = 16#11D6# else
		x"F051" when address_in = 16#11D7# else
		x"2FDB" when address_in = 16#11D8# else
		x"2FCA" when address_in = 16#11D9# else
		x"8988" when address_in = 16#11DA# else
		x"8999" when address_in = 16#11DB# else
		x"8395" when address_in = 16#11DC# else
		x"8384" when address_in = 16#11DD# else
		x"8183" when address_in = 16#11DE# else
		x"5081" when address_in = 16#11DF# else
		x"8383" when address_in = 16#11E0# else
		x"C020" when address_in = 16#11E1# else
		x"85A0" when address_in = 16#11E2# else
		x"85B1" when address_in = 16#11E3# else
		x"9710" when address_in = 16#11E4# else
		x"F051" when address_in = 16#11E5# else
		x"2FDB" when address_in = 16#11E6# else
		x"2FCA" when address_in = 16#11E7# else
		x"8988" when address_in = 16#11E8# else
		x"8999" when address_in = 16#11E9# else
		x"8791" when address_in = 16#11EA# else
		x"8780" when address_in = 16#11EB# else
		x"8182" when address_in = 16#11EC# else
		x"5081" when address_in = 16#11ED# else
		x"8382" when address_in = 16#11EE# else
		x"C012" when address_in = 16#11EF# else
		x"85A4" when address_in = 16#11F0# else
		x"85B5" when address_in = 16#11F1# else
		x"9710" when address_in = 16#11F2# else
		x"F051" when address_in = 16#11F3# else
		x"2FDB" when address_in = 16#11F4# else
		x"2FCA" when address_in = 16#11F5# else
		x"8988" when address_in = 16#11F6# else
		x"8999" when address_in = 16#11F7# else
		x"8795" when address_in = 16#11F8# else
		x"8784" when address_in = 16#11F9# else
		x"8181" when address_in = 16#11FA# else
		x"5081" when address_in = 16#11FB# else
		x"8381" when address_in = 16#11FC# else
		x"C004" when address_in = 16#11FD# else
		x"BF2F" when address_in = 16#11FE# else
		x"E080" when address_in = 16#11FF# else
		x"E090" when address_in = 16#1200# else
		x"C006" when address_in = 16#1201# else
		x"8180" when address_in = 16#1202# else
		x"5081" when address_in = 16#1203# else
		x"8380" when address_in = 16#1204# else
		x"BF2F" when address_in = 16#1205# else
		x"2F8A" when address_in = 16#1206# else
		x"2F9B" when address_in = 16#1207# else
		x"91DF" when address_in = 16#1208# else
		x"91CF" when address_in = 16#1209# else
		x"9508" when address_in = 16#120A# else
		x"92AF" when address_in = 16#120B# else
		x"92BF" when address_in = 16#120C# else
		x"92CF" when address_in = 16#120D# else
		x"92DF" when address_in = 16#120E# else
		x"92EF" when address_in = 16#120F# else
		x"92FF" when address_in = 16#1210# else
		x"930F" when address_in = 16#1211# else
		x"931F" when address_in = 16#1212# else
		x"93CF" when address_in = 16#1213# else
		x"93DF" when address_in = 16#1214# else
		x"2EE8" when address_in = 16#1215# else
		x"2EF9" when address_in = 16#1216# else
		x"2F06" when address_in = 16#1217# else
		x"2F17" when address_in = 16#1218# else
		x"2FB5" when address_in = 16#1219# else
		x"2FA4" when address_in = 16#121A# else
		x"2FD9" when address_in = 16#121B# else
		x"2FC8" when address_in = 16#121C# else
		x"81E8" when address_in = 16#121D# else
		x"81F9" when address_in = 16#121E# else
		x"2ECE" when address_in = 16#121F# else
		x"2EDF" when address_in = 16#1220# else
		x"2F6E" when address_in = 16#1221# else
		x"2F7F" when address_in = 16#1222# else
		x"9730" when address_in = 16#1223# else
		x"F409" when address_in = 16#1224# else
		x"C069" when address_in = 16#1225# else
		x"919C" when address_in = 16#1226# else
		x"8180" when address_in = 16#1227# else
		x"1798" when address_in = 16#1228# else
		x"F009" when address_in = 16#1229# else
		x"C05E" when address_in = 16#122A# else
		x"2FDB" when address_in = 16#122B# else
		x"2FCA" when address_in = 16#122C# else
		x"8199" when address_in = 16#122D# else
		x"8181" when address_in = 16#122E# else
		x"1798" when address_in = 16#122F# else
		x"F009" when address_in = 16#1230# else
		x"C057" when address_in = 16#1231# else
		x"812A" when address_in = 16#1232# else
		x"813B" when address_in = 16#1233# else
		x"8182" when address_in = 16#1234# else
		x"8193" when address_in = 16#1235# else
		x"1728" when address_in = 16#1236# else
		x"0739" when address_in = 16#1237# else
		x"F009" when address_in = 16#1238# else
		x"C04F" when address_in = 16#1239# else
		x"812C" when address_in = 16#123A# else
		x"813D" when address_in = 16#123B# else
		x"8184" when address_in = 16#123C# else
		x"8195" when address_in = 16#123D# else
		x"1728" when address_in = 16#123E# else
		x"0739" when address_in = 16#123F# else
		x"F009" when address_in = 16#1240# else
		x"C047" when address_in = 16#1241# else
		x"819E" when address_in = 16#1242# else
		x"8186" when address_in = 16#1243# else
		x"1798" when address_in = 16#1244# else
		x"F009" when address_in = 16#1245# else
		x"C042" when address_in = 16#1246# else
		x"814F" when address_in = 16#1247# else
		x"8187" when address_in = 16#1248# else
		x"1748" when address_in = 16#1249# else
		x"F5F1" when address_in = 16#124A# else
		x"E050" when address_in = 16#124B# else
		x"1754" when address_in = 16#124C# else
		x"F498" when address_in = 16#124D# else
		x"8520" when address_in = 16#124E# else
		x"8531" when address_in = 16#124F# else
		x"84A8" when address_in = 16#1250# else
		x"84B9" when address_in = 16#1251# else
		x"2DDB" when address_in = 16#1252# else
		x"2DCA" when address_in = 16#1253# else
		x"9199" when address_in = 16#1254# else
		x"2EAC" when address_in = 16#1255# else
		x"2EBD" when address_in = 16#1256# else
		x"2FD3" when address_in = 16#1257# else
		x"2FC2" when address_in = 16#1258# else
		x"9189" when address_in = 16#1259# else
		x"2F2C" when address_in = 16#125A# else
		x"2F3D" when address_in = 16#125B# else
		x"1798" when address_in = 16#125C# else
		x"F559" when address_in = 16#125D# else
		x"5F5F" when address_in = 16#125E# else
		x"1754" when address_in = 16#125F# else
		x"F388" when address_in = 16#1260# else
		x"15EC" when address_in = 16#1261# else
		x"05FD" when address_in = 16#1262# else
		x"F469" when address_in = 16#1263# else
		x"8980" when address_in = 16#1264# else
		x"8991" when address_in = 16#1265# else
		x"2DBF" when address_in = 16#1266# else
		x"2DAE" when address_in = 16#1267# else
		x"938D" when address_in = 16#1268# else
		x"939C" when address_in = 16#1269# else
		x"9700" when address_in = 16#126A# else
		x"F4D1" when address_in = 16#126B# else
		x"2FD1" when address_in = 16#126C# else
		x"2FC0" when address_in = 16#126D# else
		x"8399" when address_in = 16#126E# else
		x"8388" when address_in = 16#126F# else
		x"C015" when address_in = 16#1270# else
		x"2FB1" when address_in = 16#1271# else
		x"2FA0" when address_in = 16#1272# else
		x"918D" when address_in = 16#1273# else
		x"919C" when address_in = 16#1274# else
		x"9711" when address_in = 16#1275# else
		x"17E8" when address_in = 16#1276# else
		x"07F9" when address_in = 16#1277# else
		x"F439" when address_in = 16#1278# else
		x"2FD7" when address_in = 16#1279# else
		x"2FC6" when address_in = 16#127A# else
		x"8A19" when address_in = 16#127B# else
		x"8A18" when address_in = 16#127C# else
		x"936D" when address_in = 16#127D# else
		x"937C" when address_in = 16#127E# else
		x"C006" when address_in = 16#127F# else
		x"8980" when address_in = 16#1280# else
		x"8991" when address_in = 16#1281# else
		x"2FD7" when address_in = 16#1282# else
		x"2FC6" when address_in = 16#1283# else
		x"8B99" when address_in = 16#1284# else
		x"8B88" when address_in = 16#1285# else
		x"2F8E" when address_in = 16#1286# else
		x"2F9F" when address_in = 16#1287# else
		x"C008" when address_in = 16#1288# else
		x"2F6E" when address_in = 16#1289# else
		x"2F7F" when address_in = 16#128A# else
		x"8800" when address_in = 16#128B# else
		x"89F1" when address_in = 16#128C# else
		x"2DE0" when address_in = 16#128D# else
		x"CF94" when address_in = 16#128E# else
		x"E080" when address_in = 16#128F# else
		x"E090" when address_in = 16#1290# else
		x"91DF" when address_in = 16#1291# else
		x"91CF" when address_in = 16#1292# else
		x"911F" when address_in = 16#1293# else
		x"910F" when address_in = 16#1294# else
		x"90FF" when address_in = 16#1295# else
		x"90EF" when address_in = 16#1296# else
		x"90DF" when address_in = 16#1297# else
		x"90CF" when address_in = 16#1298# else
		x"90BF" when address_in = 16#1299# else
		x"90AF" when address_in = 16#129A# else
		x"9508" when address_in = 16#129B# else
		x"92FF" when address_in = 16#129C# else
		x"930F" when address_in = 16#129D# else
		x"931F" when address_in = 16#129E# else
		x"93CF" when address_in = 16#129F# else
		x"93DF" when address_in = 16#12A0# else
		x"2FD9" when address_in = 16#12A1# else
		x"2FC8" when address_in = 16#12A2# else
		x"2F06" when address_in = 16#12A3# else
		x"2F17" when address_in = 16#12A4# else
		x"8188" when address_in = 16#12A5# else
		x"2388" when address_in = 16#12A6# else
		x"F419" when address_in = 16#12A7# else
		x"E080" when address_in = 16#12A8# else
		x"E090" when address_in = 16#12A9# else
		x"C02D" when address_in = 16#12AA# else
		x"B6FF" when address_in = 16#12AB# else
		x"94F8" when address_in = 16#12AC# else
		x"2F8C" when address_in = 16#12AD# else
		x"2F9D" when address_in = 16#12AE# else
		x"9606" when address_in = 16#12AF# else
		x"2F46" when address_in = 16#12B0# else
		x"2F57" when address_in = 16#12B1# else
		x"2F68" when address_in = 16#12B2# else
		x"2F79" when address_in = 16#12B3# else
		x"2F8C" when address_in = 16#12B4# else
		x"2F9D" when address_in = 16#12B5# else
		x"9604" when address_in = 16#12B6# else
		x"940E" when address_in = 16#12B7# else
		x"120B" when address_in = 16#12B8# else
		x"2F28" when address_in = 16#12B9# else
		x"2F39" when address_in = 16#12BA# else
		x"2B89" when address_in = 16#12BB# else
		x"F029" when address_in = 16#12BC# else
		x"8188" when address_in = 16#12BD# else
		x"5081" when address_in = 16#12BE# else
		x"8388" when address_in = 16#12BF# else
		x"BEFF" when address_in = 16#12C0# else
		x"C014" when address_in = 16#12C1# else
		x"2F8C" when address_in = 16#12C2# else
		x"2F9D" when address_in = 16#12C3# else
		x"960E" when address_in = 16#12C4# else
		x"2F51" when address_in = 16#12C5# else
		x"2F40" when address_in = 16#12C6# else
		x"2F68" when address_in = 16#12C7# else
		x"2F79" when address_in = 16#12C8# else
		x"2F8C" when address_in = 16#12C9# else
		x"2F9D" when address_in = 16#12CA# else
		x"960C" when address_in = 16#12CB# else
		x"940E" when address_in = 16#12CC# else
		x"120B" when address_in = 16#12CD# else
		x"2F28" when address_in = 16#12CE# else
		x"2F39" when address_in = 16#12CF# else
		x"2B89" when address_in = 16#12D0# else
		x"F019" when address_in = 16#12D1# else
		x"8188" when address_in = 16#12D2# else
		x"5081" when address_in = 16#12D3# else
		x"8388" when address_in = 16#12D4# else
		x"BEFF" when address_in = 16#12D5# else
		x"2F93" when address_in = 16#12D6# else
		x"2F82" when address_in = 16#12D7# else
		x"91DF" when address_in = 16#12D8# else
		x"91CF" when address_in = 16#12D9# else
		x"911F" when address_in = 16#12DA# else
		x"910F" when address_in = 16#12DB# else
		x"90FF" when address_in = 16#12DC# else
		x"9508" when address_in = 16#12DD# else
		x"931F" when address_in = 16#12DE# else
		x"93CF" when address_in = 16#12DF# else
		x"93DF" when address_in = 16#12E0# else
		x"E0A0" when address_in = 16#12E1# else
		x"E0B0" when address_in = 16#12E2# else
		x"2FDB" when address_in = 16#12E3# else
		x"2FCA" when address_in = 16#12E4# else
		x"B71F" when address_in = 16#12E5# else
		x"94F8" when address_in = 16#12E6# else
		x"EBE7" when address_in = 16#12E7# else
		x"E0F0" when address_in = 16#12E8# else
		x"5BE6" when address_in = 16#12E9# else
		x"4FFF" when address_in = 16#12EA# else
		x"8180" when address_in = 16#12EB# else
		x"54EA" when address_in = 16#12EC# else
		x"40F0" when address_in = 16#12ED# else
		x"308F" when address_in = 16#12EE# else
		x"F439" when address_in = 16#12EF# else
		x"2FCE" when address_in = 16#12F0# else
		x"2FDF" when address_in = 16#12F1# else
		x"9001" when address_in = 16#12F2# else
		x"81F0" when address_in = 16#12F3# else
		x"2DE0" when address_in = 16#12F4# else
		x"9730" when address_in = 16#12F5# else
		x"F791" when address_in = 16#12F6# else
		x"9730" when address_in = 16#12F7# else
		x"F5B1" when address_in = 16#12F8# else
		x"B184" when address_in = 16#12F9# else
		x"2799" when address_in = 16#12FA# else
		x"718E" when address_in = 16#12FB# else
		x"7090" when address_in = 16#12FC# else
		x"9595" when address_in = 16#12FD# else
		x"9587" when address_in = 16#12FE# else
		x"9595" when address_in = 16#12FF# else
		x"9587" when address_in = 16#1300# else
		x"2F48" when address_in = 16#1301# else
		x"E06B" when address_in = 16#1302# else
		x"E48B" when address_in = 16#1303# else
		x"E090" when address_in = 16#1304# else
		x"940E" when address_in = 16#1305# else
		x"0889" when address_in = 16#1306# else
		x"8399" when address_in = 16#1307# else
		x"8388" when address_in = 16#1308# else
		x"9700" when address_in = 16#1309# else
		x"F421" when address_in = 16#130A# else
		x"BF1F" when address_in = 16#130B# else
		x"E080" when address_in = 16#130C# else
		x"E090" when address_in = 16#130D# else
		x"C03A" when address_in = 16#130E# else
		x"2FF9" when address_in = 16#130F# else
		x"2FE8" when address_in = 16#1310# else
		x"8211" when address_in = 16#1311# else
		x"8210" when address_in = 16#1312# else
		x"5BE6" when address_in = 16#1313# else
		x"4FFF" when address_in = 16#1314# else
		x"E081" when address_in = 16#1315# else
		x"8380" when address_in = 16#1316# else
		x"2FAE" when address_in = 16#1317# else
		x"2FBF" when address_in = 16#1318# else
		x"54A8" when address_in = 16#1319# else
		x"40B0" when address_in = 16#131A# else
		x"C021" when address_in = 16#131B# else
		x"2B23" when address_in = 16#131C# else
		x"8328" when address_in = 16#131D# else
		x"2F89" when address_in = 16#131E# else
		x"2799" when address_in = 16#131F# else
		x"2FB9" when address_in = 16#1320# else
		x"2FA8" when address_in = 16#1321# else
		x"E024" when address_in = 16#1322# else
		x"0FAA" when address_in = 16#1323# else
		x"1FBB" when address_in = 16#1324# else
		x"952A" when address_in = 16#1325# else
		x"F7E1" when address_in = 16#1326# else
		x"0FA8" when address_in = 16#1327# else
		x"1FB9" when address_in = 16#1328# else
		x"0FA8" when address_in = 16#1329# else
		x"1FB9" when address_in = 16#132A# else
		x"0FAE" when address_in = 16#132B# else
		x"1FBF" when address_in = 16#132C# else
		x"9612" when address_in = 16#132D# else
		x"C00E" when address_in = 16#132E# else
		x"E090" when address_in = 16#132F# else
		x"E031" when address_in = 16#1330# else
		x"2FCE" when address_in = 16#1331# else
		x"2FDF" when address_in = 16#1332# else
		x"5BC6" when address_in = 16#1333# else
		x"4FDF" when address_in = 16#1334# else
		x"8128" when address_in = 16#1335# else
		x"2F82" when address_in = 16#1336# else
		x"2383" when address_in = 16#1337# else
		x"F319" when address_in = 16#1338# else
		x"5F9F" when address_in = 16#1339# else
		x"0F33" when address_in = 16#133A# else
		x"3094" when address_in = 16#133B# else
		x"F3C8" when address_in = 16#133C# else
		x"BF1F" when address_in = 16#133D# else
		x"2F8A" when address_in = 16#133E# else
		x"2F9B" when address_in = 16#133F# else
		x"960C" when address_in = 16#1340# else
		x"2FFB" when address_in = 16#1341# else
		x"2FEA" when address_in = 16#1342# else
		x"8791" when address_in = 16#1343# else
		x"8780" when address_in = 16#1344# else
		x"8613" when address_in = 16#1345# else
		x"8612" when address_in = 16#1346# else
		x"2F8A" when address_in = 16#1347# else
		x"2F9B" when address_in = 16#1348# else
		x"91DF" when address_in = 16#1349# else
		x"91CF" when address_in = 16#134A# else
		x"911F" when address_in = 16#134B# else
		x"9508" when address_in = 16#134C# else
		x"92EF" when address_in = 16#134D# else
		x"92FF" when address_in = 16#134E# else
		x"931F" when address_in = 16#134F# else
		x"93CF" when address_in = 16#1350# else
		x"93DF" when address_in = 16#1351# else
		x"2FD9" when address_in = 16#1352# else
		x"2FC8" when address_in = 16#1353# else
		x"24EE" when address_in = 16#1354# else
		x"24FF" when address_in = 16#1355# else
		x"858A" when address_in = 16#1356# else
		x"859B" when address_in = 16#1357# else
		x"FF82" when address_in = 16#1358# else
		x"C00D" when address_in = 16#1359# else
		x"B184" when address_in = 16#135A# else
		x"2799" when address_in = 16#135B# else
		x"718E" when address_in = 16#135C# else
		x"7090" when address_in = 16#135D# else
		x"9595" when address_in = 16#135E# else
		x"9587" when address_in = 16#135F# else
		x"9595" when address_in = 16#1360# else
		x"9587" when address_in = 16#1361# else
		x"2F68" when address_in = 16#1362# else
		x"8588" when address_in = 16#1363# else
		x"8599" when address_in = 16#1364# else
		x"940E" when address_in = 16#1365# else
		x"07EC" when address_in = 16#1366# else
		x"B71F" when address_in = 16#1367# else
		x"94F8" when address_in = 16#1368# else
		x"EBA7" when address_in = 16#1369# else
		x"E0B0" when address_in = 16#136A# else
		x"2F8A" when address_in = 16#136B# else
		x"2F9B" when address_in = 16#136C# else
		x"9602" when address_in = 16#136D# else
		x"17C8" when address_in = 16#136E# else
		x"07D9" when address_in = 16#136F# else
		x"F1B8" when address_in = 16#1370# else
		x"2FFB" when address_in = 16#1371# else
		x"2FEA" when address_in = 16#1372# else
		x"5BE6" when address_in = 16#1373# else
		x"4FFF" when address_in = 16#1374# else
		x"17CE" when address_in = 16#1375# else
		x"07DF" when address_in = 16#1376# else
		x"F580" when address_in = 16#1377# else
		x"1BCA" when address_in = 16#1378# else
		x"0BDB" when address_in = 16#1379# else
		x"9722" when address_in = 16#137A# else
		x"2F8C" when address_in = 16#137B# else
		x"2F9D" when address_in = 16#137C# else
		x"9595" when address_in = 16#137D# else
		x"9587" when address_in = 16#137E# else
		x"E369" when address_in = 16#137F# else
		x"E87E" when address_in = 16#1380# else
		x"940E" when address_in = 16#1381# else
		x"2E76" when address_in = 16#1382# else
		x"E021" when address_in = 16#1383# else
		x"E030" when address_in = 16#1384# else
		x"C002" when address_in = 16#1385# else
		x"0F22" when address_in = 16#1386# else
		x"1F33" when address_in = 16#1387# else
		x"958A" when address_in = 16#1388# else
		x"F7E2" when address_in = 16#1389# else
		x"2F92" when address_in = 16#138A# else
		x"9590" when address_in = 16#138B# else
		x"8180" when address_in = 16#138C# else
		x"2389" when address_in = 16#138D# else
		x"8380" when address_in = 16#138E# else
		x"2388" when address_in = 16#138F# else
		x"F4A9" when address_in = 16#1390# else
		x"E080" when address_in = 16#1391# else
		x"3BA7" when address_in = 16#1392# else
		x"07B8" when address_in = 16#1393# else
		x"F089" when address_in = 16#1394# else
		x"B184" when address_in = 16#1395# else
		x"2799" when address_in = 16#1396# else
		x"718E" when address_in = 16#1397# else
		x"7090" when address_in = 16#1398# else
		x"9595" when address_in = 16#1399# else
		x"9587" when address_in = 16#139A# else
		x"9595" when address_in = 16#139B# else
		x"9587" when address_in = 16#139C# else
		x"2F68" when address_in = 16#139D# else
		x"2F8A" when address_in = 16#139E# else
		x"2F9B" when address_in = 16#139F# else
		x"940E" when address_in = 16#13A0# else
		x"07EC" when address_in = 16#13A1# else
		x"2DFF" when address_in = 16#13A2# else
		x"2DEE" when address_in = 16#13A3# else
		x"8211" when address_in = 16#13A4# else
		x"8210" when address_in = 16#13A5# else
		x"BF1F" when address_in = 16#13A6# else
		x"C016" when address_in = 16#13A7# else
		x"2EEA" when address_in = 16#13A8# else
		x"2EFB" when address_in = 16#13A9# else
		x"900D" when address_in = 16#13AA# else
		x"91BC" when address_in = 16#13AB# else
		x"2DA0" when address_in = 16#13AC# else
		x"9710" when address_in = 16#13AD# else
		x"F009" when address_in = 16#13AE# else
		x"CFBB" when address_in = 16#13AF# else
		x"B184" when address_in = 16#13B0# else
		x"2799" when address_in = 16#13B1# else
		x"718E" when address_in = 16#13B2# else
		x"7090" when address_in = 16#13B3# else
		x"9595" when address_in = 16#13B4# else
		x"9587" when address_in = 16#13B5# else
		x"9595" when address_in = 16#13B6# else
		x"9587" when address_in = 16#13B7# else
		x"2F68" when address_in = 16#13B8# else
		x"2F8C" when address_in = 16#13B9# else
		x"2F9D" when address_in = 16#13BA# else
		x"940E" when address_in = 16#13BB# else
		x"07EC" when address_in = 16#13BC# else
		x"BF1F" when address_in = 16#13BD# else
		x"91DF" when address_in = 16#13BE# else
		x"91CF" when address_in = 16#13BF# else
		x"911F" when address_in = 16#13C0# else
		x"90FF" when address_in = 16#13C1# else
		x"90EF" when address_in = 16#13C2# else
		x"9508" when address_in = 16#13C3# else
		x"92DF" when address_in = 16#13C4# else
		x"92EF" when address_in = 16#13C5# else
		x"92FF" when address_in = 16#13C6# else
		x"930F" when address_in = 16#13C7# else
		x"931F" when address_in = 16#13C8# else
		x"93CF" when address_in = 16#13C9# else
		x"93DF" when address_in = 16#13CA# else
		x"2FD9" when address_in = 16#13CB# else
		x"2FC8" when address_in = 16#13CC# else
		x"2F16" when address_in = 16#13CD# else
		x"2ED4" when address_in = 16#13CE# else
		x"858A" when address_in = 16#13CF# else
		x"859B" when address_in = 16#13D0# else
		x"FF83" when address_in = 16#13D1# else
		x"C028" when address_in = 16#13D2# else
		x"FF82" when address_in = 16#13D3# else
		x"C014" when address_in = 16#13D4# else
		x"B184" when address_in = 16#13D5# else
		x"2799" when address_in = 16#13D6# else
		x"718E" when address_in = 16#13D7# else
		x"7090" when address_in = 16#13D8# else
		x"9595" when address_in = 16#13D9# else
		x"9587" when address_in = 16#13DA# else
		x"9595" when address_in = 16#13DB# else
		x"9587" when address_in = 16#13DC# else
		x"2F68" when address_in = 16#13DD# else
		x"8588" when address_in = 16#13DE# else
		x"8599" when address_in = 16#13DF# else
		x"940E" when address_in = 16#13E0# else
		x"07EC" when address_in = 16#13E1# else
		x"858A" when address_in = 16#13E2# else
		x"859B" when address_in = 16#13E3# else
		x"7F8B" when address_in = 16#13E4# else
		x"879B" when address_in = 16#13E5# else
		x"878A" when address_in = 16#13E6# else
		x"8619" when address_in = 16#13E7# else
		x"8618" when address_in = 16#13E8# else
		x"2311" when address_in = 16#13E9# else
		x"F411" when address_in = 16#13EA# else
		x"E082" when address_in = 16#13EB# else
		x"C001" when address_in = 16#13EC# else
		x"E080" when address_in = 16#13ED# else
		x"2799" when address_in = 16#13EE# else
		x"2EE8" when address_in = 16#13EF# else
		x"2EF9" when address_in = 16#13F0# else
		x"2F0C" when address_in = 16#13F1# else
		x"2F1D" when address_in = 16#13F2# else
		x"E122" when address_in = 16#13F3# else
		x"E043" when address_in = 16#13F4# else
		x"2D6D" when address_in = 16#13F5# else
		x"8189" when address_in = 16#13F6# else
		x"940E" when address_in = 16#13F7# else
		x"105C" when address_in = 16#13F8# else
		x"FF87" when address_in = 16#13F9# else
		x"C004" when address_in = 16#13FA# else
		x"2F8C" when address_in = 16#13FB# else
		x"2F9D" when address_in = 16#13FC# else
		x"940E" when address_in = 16#13FD# else
		x"134D" when address_in = 16#13FE# else
		x"91DF" when address_in = 16#13FF# else
		x"91CF" when address_in = 16#1400# else
		x"911F" when address_in = 16#1401# else
		x"910F" when address_in = 16#1402# else
		x"90FF" when address_in = 16#1403# else
		x"90EF" when address_in = 16#1404# else
		x"90DF" when address_in = 16#1405# else
		x"9508" when address_in = 16#1406# else
		x"92FF" when address_in = 16#1407# else
		x"930F" when address_in = 16#1408# else
		x"931F" when address_in = 16#1409# else
		x"93CF" when address_in = 16#140A# else
		x"93DF" when address_in = 16#140B# else
		x"B7CD" when address_in = 16#140C# else
		x"B7DE" when address_in = 16#140D# else
		x"9728" when address_in = 16#140E# else
		x"B60F" when address_in = 16#140F# else
		x"94F8" when address_in = 16#1410# else
		x"BFDE" when address_in = 16#1411# else
		x"BE0F" when address_in = 16#1412# else
		x"BFCD" when address_in = 16#1413# else
		x"2F08" when address_in = 16#1414# else
		x"2F19" when address_in = 16#1415# else
		x"E088" when address_in = 16#1416# else
		x"2FFD" when address_in = 16#1417# else
		x"2FEC" when address_in = 16#1418# else
		x"9631" when address_in = 16#1419# else
		x"9211" when address_in = 16#141A# else
		x"958A" when address_in = 16#141B# else
		x"F7E9" when address_in = 16#141C# else
		x"9180" when address_in = 16#141D# else
		x"0062" when address_in = 16#141E# else
		x"9190" when address_in = 16#141F# else
		x"0063" when address_in = 16#1420# else
		x"2FF1" when address_in = 16#1421# else
		x"2FE0" when address_in = 16#1422# else
		x"8122" when address_in = 16#1423# else
		x"8133" when address_in = 16#1424# else
		x"1782" when address_in = 16#1425# else
		x"0793" when address_in = 16#1426# else
		x"F429" when address_in = 16#1427# else
		x"2F91" when address_in = 16#1428# else
		x"2F80" when address_in = 16#1429# else
		x"940E" when address_in = 16#142A# else
		x"0EC0" when address_in = 16#142B# else
		x"C051" when address_in = 16#142C# else
		x"2FF1" when address_in = 16#142D# else
		x"2FE0" when address_in = 16#142E# else
		x"8582" when address_in = 16#142F# else
		x"8593" when address_in = 16#1430# else
		x"FF95" when address_in = 16#1431# else
		x"C02E" when address_in = 16#1432# else
		x"EFFF" when address_in = 16#1433# else
		x"3F2F" when address_in = 16#1434# else
		x"073F" when address_in = 16#1435# else
		x"F151" when address_in = 16#1436# else
		x"24FF" when address_in = 16#1437# else
		x"2F93" when address_in = 16#1438# else
		x"2F82" when address_in = 16#1439# else
		x"940E" when address_in = 16#143A# else
		x"26BD" when address_in = 16#143B# else
		x"2FF1" when address_in = 16#143C# else
		x"2FE0" when address_in = 16#143D# else
		x"8522" when address_in = 16#143E# else
		x"8533" when address_in = 16#143F# else
		x"2388" when address_in = 16#1440# else
		x"F431" when address_in = 16#1441# else
		x"6038" when address_in = 16#1442# else
		x"8733" when address_in = 16#1443# else
		x"8722" when address_in = 16#1444# else
		x"E081" when address_in = 16#1445# else
		x"2EF8" when address_in = 16#1446# else
		x"C005" when address_in = 16#1447# else
		x"7F37" when address_in = 16#1448# else
		x"2FF1" when address_in = 16#1449# else
		x"2FE0" when address_in = 16#144A# else
		x"8733" when address_in = 16#144B# else
		x"8722" when address_in = 16#144C# else
		x"2FF1" when address_in = 16#144D# else
		x"2FE0" when address_in = 16#144E# else
		x"8522" when address_in = 16#144F# else
		x"8533" when address_in = 16#1450# else
		x"2F93" when address_in = 16#1451# else
		x"2F82" when address_in = 16#1452# else
		x"7F9B" when address_in = 16#1453# else
		x"8793" when address_in = 16#1454# else
		x"8782" when address_in = 16#1455# else
		x"20FF" when address_in = 16#1456# else
		x"F421" when address_in = 16#1457# else
		x"6092" when address_in = 16#1458# else
		x"8793" when address_in = 16#1459# else
		x"8782" when address_in = 16#145A# else
		x"C005" when address_in = 16#145B# else
		x"7F39" when address_in = 16#145C# else
		x"2FF1" when address_in = 16#145D# else
		x"2FE0" when address_in = 16#145E# else
		x"8733" when address_in = 16#145F# else
		x"8722" when address_in = 16#1460# else
		x"2FF1" when address_in = 16#1461# else
		x"2FE0" when address_in = 16#1462# else
		x"8522" when address_in = 16#1463# else
		x"8533" when address_in = 16#1464# else
		x"2F93" when address_in = 16#1465# else
		x"2F82" when address_in = 16#1466# else
		x"7080" when address_in = 16#1467# else
		x"719E" when address_in = 16#1468# else
		x"2B89" when address_in = 16#1469# else
		x"F429" when address_in = 16#146A# else
		x"2F91" when address_in = 16#146B# else
		x"2F80" when address_in = 16#146C# else
		x"940E" when address_in = 16#146D# else
		x"134D" when address_in = 16#146E# else
		x"C00E" when address_in = 16#146F# else
		x"FF33" when address_in = 16#1470# else
		x"C002" when address_in = 16#1471# else
		x"831E" when address_in = 16#1472# else
		x"830D" when address_in = 16#1473# else
		x"2F91" when address_in = 16#1474# else
		x"2F80" when address_in = 16#1475# else
		x"940E" when address_in = 16#1476# else
		x"236F" when address_in = 16#1477# else
		x"818D" when address_in = 16#1478# else
		x"819E" when address_in = 16#1479# else
		x"9700" when address_in = 16#147A# else
		x"F011" when address_in = 16#147B# else
		x"940E" when address_in = 16#147C# else
		x"25F8" when address_in = 16#147D# else
		x"E080" when address_in = 16#147E# else
		x"E090" when address_in = 16#147F# else
		x"9628" when address_in = 16#1480# else
		x"B60F" when address_in = 16#1481# else
		x"94F8" when address_in = 16#1482# else
		x"BFDE" when address_in = 16#1483# else
		x"BE0F" when address_in = 16#1484# else
		x"BFCD" when address_in = 16#1485# else
		x"91DF" when address_in = 16#1486# else
		x"91CF" when address_in = 16#1487# else
		x"911F" when address_in = 16#1488# else
		x"910F" when address_in = 16#1489# else
		x"90FF" when address_in = 16#148A# else
		x"9508" when address_in = 16#148B# else
		x"929F" when address_in = 16#148C# else
		x"92AF" when address_in = 16#148D# else
		x"92BF" when address_in = 16#148E# else
		x"92CF" when address_in = 16#148F# else
		x"92DF" when address_in = 16#1490# else
		x"92EF" when address_in = 16#1491# else
		x"92FF" when address_in = 16#1492# else
		x"930F" when address_in = 16#1493# else
		x"931F" when address_in = 16#1494# else
		x"93CF" when address_in = 16#1495# else
		x"2EB8" when address_in = 16#1496# else
		x"2E96" when address_in = 16#1497# else
		x"2FC4" when address_in = 16#1498# else
		x"2EA2" when address_in = 16#1499# else
		x"940E" when address_in = 16#149A# else
		x"12DE" when address_in = 16#149B# else
		x"2FF9" when address_in = 16#149C# else
		x"2FE8" when address_in = 16#149D# else
		x"2B89" when address_in = 16#149E# else
		x"F491" when address_in = 16#149F# else
		x"FEE2" when address_in = 16#14A0# else
		x"C00D" when address_in = 16#14A1# else
		x"B184" when address_in = 16#14A2# else
		x"2799" when address_in = 16#14A3# else
		x"718E" when address_in = 16#14A4# else
		x"7090" when address_in = 16#14A5# else
		x"9595" when address_in = 16#14A6# else
		x"9587" when address_in = 16#14A7# else
		x"9595" when address_in = 16#14A8# else
		x"9587" when address_in = 16#14A9# else
		x"2F68" when address_in = 16#14AA# else
		x"2F91" when address_in = 16#14AB# else
		x"2F80" when address_in = 16#14AC# else
		x"940E" when address_in = 16#14AD# else
		x"07EC" when address_in = 16#14AE# else
		x"EF84" when address_in = 16#14AF# else
		x"EF9F" when address_in = 16#14B0# else
		x"C017" when address_in = 16#14B1# else
		x"82D3" when address_in = 16#14B2# else
		x"82C2" when address_in = 16#14B3# else
		x"82B0" when address_in = 16#14B4# else
		x"83C6" when address_in = 16#14B5# else
		x"9180" when address_in = 16#14B6# else
		x"0062" when address_in = 16#14B7# else
		x"9190" when address_in = 16#14B8# else
		x"0063" when address_in = 16#14B9# else
		x"8395" when address_in = 16#14BA# else
		x"8384" when address_in = 16#14BB# else
		x"8291" when address_in = 16#14BC# else
		x"82A7" when address_in = 16#14BD# else
		x"8711" when address_in = 16#14BE# else
		x"8700" when address_in = 16#14BF# else
		x"86F3" when address_in = 16#14C0# else
		x"86E2" when address_in = 16#14C1# else
		x"2F8E" when address_in = 16#14C2# else
		x"2F9F" when address_in = 16#14C3# else
		x"940E" when address_in = 16#14C4# else
		x"1407" when address_in = 16#14C5# else
		x"2799" when address_in = 16#14C6# else
		x"FD87" when address_in = 16#14C7# else
		x"9590" when address_in = 16#14C8# else
		x"91CF" when address_in = 16#14C9# else
		x"911F" when address_in = 16#14CA# else
		x"910F" when address_in = 16#14CB# else
		x"90FF" when address_in = 16#14CC# else
		x"90EF" when address_in = 16#14CD# else
		x"90DF" when address_in = 16#14CE# else
		x"90CF" when address_in = 16#14CF# else
		x"90BF" when address_in = 16#14D0# else
		x"90AF" when address_in = 16#14D1# else
		x"909F" when address_in = 16#14D2# else
		x"9508" when address_in = 16#14D3# else
		x"93CF" when address_in = 16#14D4# else
		x"93DF" when address_in = 16#14D5# else
		x"2FD9" when address_in = 16#14D6# else
		x"2FC8" when address_in = 16#14D7# else
		x"940E" when address_in = 16#14D8# else
		x"12DE" when address_in = 16#14D9# else
		x"2FF9" when address_in = 16#14DA# else
		x"2FE8" when address_in = 16#14DB# else
		x"2B89" when address_in = 16#14DC# else
		x"F4A1" when address_in = 16#14DD# else
		x"858A" when address_in = 16#14DE# else
		x"859B" when address_in = 16#14DF# else
		x"FF82" when address_in = 16#14E0# else
		x"C00D" when address_in = 16#14E1# else
		x"B184" when address_in = 16#14E2# else
		x"2799" when address_in = 16#14E3# else
		x"718E" when address_in = 16#14E4# else
		x"7090" when address_in = 16#14E5# else
		x"9595" when address_in = 16#14E6# else
		x"9587" when address_in = 16#14E7# else
		x"9595" when address_in = 16#14E8# else
		x"9587" when address_in = 16#14E9# else
		x"2F68" when address_in = 16#14EA# else
		x"8588" when address_in = 16#14EB# else
		x"8599" when address_in = 16#14EC# else
		x"940E" when address_in = 16#14ED# else
		x"07EC" when address_in = 16#14EE# else
		x"EF84" when address_in = 16#14EF# else
		x"EF9F" when address_in = 16#14F0# else
		x"C00E" when address_in = 16#14F1# else
		x"E182" when address_in = 16#14F2# else
		x"2FAE" when address_in = 16#14F3# else
		x"2FBF" when address_in = 16#14F4# else
		x"9009" when address_in = 16#14F5# else
		x"920D" when address_in = 16#14F6# else
		x"958A" when address_in = 16#14F7# else
		x"F7E1" when address_in = 16#14F8# else
		x"2F8E" when address_in = 16#14F9# else
		x"2F9F" when address_in = 16#14FA# else
		x"940E" when address_in = 16#14FB# else
		x"1407" when address_in = 16#14FC# else
		x"2799" when address_in = 16#14FD# else
		x"FD87" when address_in = 16#14FE# else
		x"9590" when address_in = 16#14FF# else
		x"91DF" when address_in = 16#1500# else
		x"91CF" when address_in = 16#1501# else
		x"9508" when address_in = 16#1502# else
		x"925F" when address_in = 16#1503# else
		x"926F" when address_in = 16#1504# else
		x"927F" when address_in = 16#1505# else
		x"928F" when address_in = 16#1506# else
		x"929F" when address_in = 16#1507# else
		x"92AF" when address_in = 16#1508# else
		x"92BF" when address_in = 16#1509# else
		x"92CF" when address_in = 16#150A# else
		x"92DF" when address_in = 16#150B# else
		x"92EF" when address_in = 16#150C# else
		x"92FF" when address_in = 16#150D# else
		x"930F" when address_in = 16#150E# else
		x"931F" when address_in = 16#150F# else
		x"93CF" when address_in = 16#1510# else
		x"2E58" when address_in = 16#1511# else
		x"2E66" when address_in = 16#1512# else
		x"2E74" when address_in = 16#1513# else
		x"2E82" when address_in = 16#1514# else
		x"2E93" when address_in = 16#1515# else
		x"2EA0" when address_in = 16#1516# else
		x"2EB1" when address_in = 16#1517# else
		x"940E" when address_in = 16#1518# else
		x"0B5D" when address_in = 16#1519# else
		x"2FC8" when address_in = 16#151A# else
		x"2CCE" when address_in = 16#151B# else
		x"2CDF" when address_in = 16#151C# else
		x"2CFB" when address_in = 16#151D# else
		x"2CEA" when address_in = 16#151E# else
		x"2D19" when address_in = 16#151F# else
		x"2D08" when address_in = 16#1520# else
		x"2D27" when address_in = 16#1521# else
		x"2D46" when address_in = 16#1522# else
		x"2F68" when address_in = 16#1523# else
		x"2D85" when address_in = 16#1524# else
		x"940E" when address_in = 16#1525# else
		x"148C" when address_in = 16#1526# else
		x"2388" when address_in = 16#1527# else
		x"F039" when address_in = 16#1528# else
		x"2F8C" when address_in = 16#1529# else
		x"940E" when address_in = 16#152A# else
		x"09FA" when address_in = 16#152B# else
		x"2799" when address_in = 16#152C# else
		x"FD87" when address_in = 16#152D# else
		x"9590" when address_in = 16#152E# else
		x"C002" when address_in = 16#152F# else
		x"E080" when address_in = 16#1530# else
		x"E090" when address_in = 16#1531# else
		x"91CF" when address_in = 16#1532# else
		x"911F" when address_in = 16#1533# else
		x"910F" when address_in = 16#1534# else
		x"90FF" when address_in = 16#1535# else
		x"90EF" when address_in = 16#1536# else
		x"90DF" when address_in = 16#1537# else
		x"90CF" when address_in = 16#1538# else
		x"90BF" when address_in = 16#1539# else
		x"90AF" when address_in = 16#153A# else
		x"909F" when address_in = 16#153B# else
		x"908F" when address_in = 16#153C# else
		x"907F" when address_in = 16#153D# else
		x"906F" when address_in = 16#153E# else
		x"905F" when address_in = 16#153F# else
		x"9508" when address_in = 16#1540# else
		x"E080" when address_in = 16#1541# else
		x"E090" when address_in = 16#1542# else
		x"9508" when address_in = 16#1543# else
		x"930F" when address_in = 16#1544# else
		x"931F" when address_in = 16#1545# else
		x"93CF" when address_in = 16#1546# else
		x"2FF9" when address_in = 16#1547# else
		x"2FE8" when address_in = 16#1548# else
		x"2F06" when address_in = 16#1549# else
		x"2F84" when address_in = 16#154A# else
		x"2F12" when address_in = 16#154B# else
		x"2FC4" when address_in = 16#154C# else
		x"1742" when address_in = 16#154D# else
		x"F5B0" when address_in = 16#154E# else
		x"2F2E" when address_in = 16#154F# else
		x"2F3F" when address_in = 16#1550# else
		x"2744" when address_in = 16#1551# else
		x"2755" when address_in = 16#1552# else
		x"0F22" when address_in = 16#1553# else
		x"1F33" when address_in = 16#1554# else
		x"1F44" when address_in = 16#1555# else
		x"1F55" when address_in = 16#1556# else
		x"2F68" when address_in = 16#1557# else
		x"2777" when address_in = 16#1558# else
		x"E093" when address_in = 16#1559# else
		x"0F66" when address_in = 16#155A# else
		x"1F77" when address_in = 16#155B# else
		x"959A" when address_in = 16#155C# else
		x"F7E1" when address_in = 16#155D# else
		x"5F69" when address_in = 16#155E# else
		x"4F7F" when address_in = 16#155F# else
		x"2F86" when address_in = 16#1560# else
		x"2F97" when address_in = 16#1561# else
		x"27AA" when address_in = 16#1562# else
		x"27BB" when address_in = 16#1563# else
		x"5067" when address_in = 16#1564# else
		x"4070" when address_in = 16#1565# else
		x"0F82" when address_in = 16#1566# else
		x"1F93" when address_in = 16#1567# else
		x"1FA4" when address_in = 16#1568# else
		x"1FB5" when address_in = 16#1569# else
		x"BFAB" when address_in = 16#156A# else
		x"2FF9" when address_in = 16#156B# else
		x"2FE8" when address_in = 16#156C# else
		x"95D8" when address_in = 16#156D# else
		x"2D80" when address_in = 16#156E# else
		x"1780" when address_in = 16#156F# else
		x"F479" when address_in = 16#1570# else
		x"2F86" when address_in = 16#1571# else
		x"2F97" when address_in = 16#1572# else
		x"27AA" when address_in = 16#1573# else
		x"27BB" when address_in = 16#1574# else
		x"0F28" when address_in = 16#1575# else
		x"1F39" when address_in = 16#1576# else
		x"1F4A" when address_in = 16#1577# else
		x"1F5B" when address_in = 16#1578# else
		x"9556" when address_in = 16#1579# else
		x"9547" when address_in = 16#157A# else
		x"9537" when address_in = 16#157B# else
		x"9527" when address_in = 16#157C# else
		x"2F93" when address_in = 16#157D# else
		x"2F82" when address_in = 16#157E# else
		x"C007" when address_in = 16#157F# else
		x"5FCF" when address_in = 16#1580# else
		x"5F68" when address_in = 16#1581# else
		x"4F7F" when address_in = 16#1582# else
		x"17C1" when address_in = 16#1583# else
		x"F2C8" when address_in = 16#1584# else
		x"E080" when address_in = 16#1585# else
		x"E090" when address_in = 16#1586# else
		x"91CF" when address_in = 16#1587# else
		x"911F" when address_in = 16#1588# else
		x"910F" when address_in = 16#1589# else
		x"9508" when address_in = 16#158A# else
		x"93CF" when address_in = 16#158B# else
		x"93DF" when address_in = 16#158C# else
		x"2FF9" when address_in = 16#158D# else
		x"2FE8" when address_in = 16#158E# else
		x"2FB7" when address_in = 16#158F# else
		x"2FA6" when address_in = 16#1590# else
		x"8190" when address_in = 16#1591# else
		x"918C" when address_in = 16#1592# else
		x"1798" when address_in = 16#1593# else
		x"F489" when address_in = 16#1594# else
		x"8191" when address_in = 16#1595# else
		x"2FD7" when address_in = 16#1596# else
		x"2FC6" when address_in = 16#1597# else
		x"8189" when address_in = 16#1598# else
		x"1798" when address_in = 16#1599# else
		x"F459" when address_in = 16#159A# else
		x"8192" when address_in = 16#159B# else
		x"818A" when address_in = 16#159C# else
		x"1798" when address_in = 16#159D# else
		x"F439" when address_in = 16#159E# else
		x"8193" when address_in = 16#159F# else
		x"818B" when address_in = 16#15A0# else
		x"1798" when address_in = 16#15A1# else
		x"F419" when address_in = 16#15A2# else
		x"E081" when address_in = 16#15A3# else
		x"E090" when address_in = 16#15A4# else
		x"C002" when address_in = 16#15A5# else
		x"E080" when address_in = 16#15A6# else
		x"E090" when address_in = 16#15A7# else
		x"91DF" when address_in = 16#15A8# else
		x"91CF" when address_in = 16#15A9# else
		x"9508" when address_in = 16#15AA# else
		x"927F" when address_in = 16#15AB# else
		x"928F" when address_in = 16#15AC# else
		x"929F" when address_in = 16#15AD# else
		x"92AF" when address_in = 16#15AE# else
		x"92BF" when address_in = 16#15AF# else
		x"92CF" when address_in = 16#15B0# else
		x"92DF" when address_in = 16#15B1# else
		x"92EF" when address_in = 16#15B2# else
		x"92FF" when address_in = 16#15B3# else
		x"930F" when address_in = 16#15B4# else
		x"931F" when address_in = 16#15B5# else
		x"93CF" when address_in = 16#15B6# else
		x"93DF" when address_in = 16#15B7# else
		x"B7CD" when address_in = 16#15B8# else
		x"B7DE" when address_in = 16#15B9# else
		x"9728" when address_in = 16#15BA# else
		x"B60F" when address_in = 16#15BB# else
		x"94F8" when address_in = 16#15BC# else
		x"BFDE" when address_in = 16#15BD# else
		x"BE0F" when address_in = 16#15BE# else
		x"BFCD" when address_in = 16#15BF# else
		x"2EC8" when address_in = 16#15C0# else
		x"2ED9" when address_in = 16#15C1# else
		x"2F86" when address_in = 16#15C2# else
		x"2F14" when address_in = 16#15C3# else
		x"2EB2" when address_in = 16#15C4# else
		x"2488" when address_in = 16#15C5# else
		x"2499" when address_in = 16#15C6# else
		x"2477" when address_in = 16#15C7# else
		x"940E" when address_in = 16#15C8# else
		x"0B28" when address_in = 16#15C9# else
		x"2FF9" when address_in = 16#15CA# else
		x"2FE8" when address_in = 16#15CB# else
		x"2B89" when address_in = 16#15CC# else
		x"F409" when address_in = 16#15CD# else
		x"C084" when address_in = 16#15CE# else
		x"8182" when address_in = 16#15CF# else
		x"8193" when address_in = 16#15D0# else
		x"27AA" when address_in = 16#15D1# else
		x"27BB" when address_in = 16#15D2# else
		x"0F88" when address_in = 16#15D3# else
		x"1F99" when address_in = 16#15D4# else
		x"1FAA" when address_in = 16#15D5# else
		x"1FBB" when address_in = 16#15D6# else
		x"9603" when address_in = 16#15D7# else
		x"1DA1" when address_in = 16#15D8# else
		x"1DB1" when address_in = 16#15D9# else
		x"BFAB" when address_in = 16#15DA# else
		x"2FF9" when address_in = 16#15DB# else
		x"2FE8" when address_in = 16#15DC# else
		x"95D8" when address_in = 16#15DD# else
		x"2D30" when address_in = 16#15DE# else
		x"9601" when address_in = 16#15DF# else
		x"1DA1" when address_in = 16#15E0# else
		x"1DB1" when address_in = 16#15E1# else
		x"BFAB" when address_in = 16#15E2# else
		x"2FF9" when address_in = 16#15E3# else
		x"2FE8" when address_in = 16#15E4# else
		x"95D8" when address_in = 16#15E5# else
		x"2D20" when address_in = 16#15E6# else
		x"0F23" when address_in = 16#15E7# else
		x"960A" when address_in = 16#15E8# else
		x"1DA1" when address_in = 16#15E9# else
		x"1DB1" when address_in = 16#15EA# else
		x"95B6" when address_in = 16#15EB# else
		x"95A7" when address_in = 16#15EC# else
		x"9597" when address_in = 16#15ED# else
		x"9587" when address_in = 16#15EE# else
		x"2F43" when address_in = 16#15EF# else
		x"2F61" when address_in = 16#15F0# else
		x"940E" when address_in = 16#15F1# else
		x"1544" when address_in = 16#15F2# else
		x"2E88" when address_in = 16#15F3# else
		x"2E99" when address_in = 16#15F4# else
		x"9700" when address_in = 16#15F5# else
		x"F409" when address_in = 16#15F6# else
		x"C05B" when address_in = 16#15F7# else
		x"2EE8" when address_in = 16#15F8# else
		x"2EF9" when address_in = 16#15F9# else
		x"2700" when address_in = 16#15FA# else
		x"2711" when address_in = 16#15FB# else
		x"0CEE" when address_in = 16#15FC# else
		x"1CFF" when address_in = 16#15FD# else
		x"1F00" when address_in = 16#15FE# else
		x"1F11" when address_in = 16#15FF# else
		x"2D4C" when address_in = 16#1600# else
		x"2D5D" when address_in = 16#1601# else
		x"2766" when address_in = 16#1602# else
		x"2777" when address_in = 16#1603# else
		x"0F44" when address_in = 16#1604# else
		x"1F55" when address_in = 16#1605# else
		x"1F66" when address_in = 16#1606# else
		x"1F77" when address_in = 16#1607# else
		x"2D2B" when address_in = 16#1608# else
		x"2733" when address_in = 16#1609# else
		x"E0E3" when address_in = 16#160A# else
		x"0F22" when address_in = 16#160B# else
		x"1F33" when address_in = 16#160C# else
		x"95EA" when address_in = 16#160D# else
		x"F7E1" when address_in = 16#160E# else
		x"5F20" when address_in = 16#160F# else
		x"4F3F" when address_in = 16#1610# else
		x"2EAC" when address_in = 16#1611# else
		x"2EBD" when address_in = 16#1612# else
		x"9408" when address_in = 16#1613# else
		x"1CA1" when address_in = 16#1614# else
		x"1CB1" when address_in = 16#1615# else
		x"24CC" when address_in = 16#1616# else
		x"24DD" when address_in = 16#1617# else
		x"E082" when address_in = 16#1618# else
		x"E090" when address_in = 16#1619# else
		x"0EC8" when address_in = 16#161A# else
		x"1ED9" when address_in = 16#161B# else
		x"2D8C" when address_in = 16#161C# else
		x"2D9D" when address_in = 16#161D# else
		x"27AA" when address_in = 16#161E# else
		x"27BB" when address_in = 16#161F# else
		x"0D8E" when address_in = 16#1620# else
		x"1D9F" when address_in = 16#1621# else
		x"1FA0" when address_in = 16#1622# else
		x"1FB1" when address_in = 16#1623# else
		x"BFAB" when address_in = 16#1624# else
		x"2FF9" when address_in = 16#1625# else
		x"2FE8" when address_in = 16#1626# else
		x"95D8" when address_in = 16#1627# else
		x"2D80" when address_in = 16#1628# else
		x"2DFB" when address_in = 16#1629# else
		x"2DEA" when address_in = 16#162A# else
		x"8380" when address_in = 16#162B# else
		x"2F82" when address_in = 16#162C# else
		x"2F93" when address_in = 16#162D# else
		x"27AA" when address_in = 16#162E# else
		x"27BB" when address_in = 16#162F# else
		x"0F84" when address_in = 16#1630# else
		x"1F95" when address_in = 16#1631# else
		x"1FA6" when address_in = 16#1632# else
		x"1FB7" when address_in = 16#1633# else
		x"BFAB" when address_in = 16#1634# else
		x"2FF9" when address_in = 16#1635# else
		x"2FE8" when address_in = 16#1636# else
		x"95D8" when address_in = 16#1637# else
		x"2D80" when address_in = 16#1638# else
		x"2DFB" when address_in = 16#1639# else
		x"2DEA" when address_in = 16#163A# else
		x"8384" when address_in = 16#163B# else
		x"9473" when address_in = 16#163C# else
		x"9408" when address_in = 16#163D# else
		x"08C1" when address_in = 16#163E# else
		x"08D1" when address_in = 16#163F# else
		x"9408" when address_in = 16#1640# else
		x"1CA1" when address_in = 16#1641# else
		x"1CB1" when address_in = 16#1642# else
		x"5F2F" when address_in = 16#1643# else
		x"4F3F" when address_in = 16#1644# else
		x"E0F3" when address_in = 16#1645# else
		x"15F7" when address_in = 16#1646# else
		x"F680" when address_in = 16#1647# else
		x"2F6C" when address_in = 16#1648# else
		x"2F7D" when address_in = 16#1649# else
		x"5F6B" when address_in = 16#164A# else
		x"4F7F" when address_in = 16#164B# else
		x"2F8C" when address_in = 16#164C# else
		x"2F9D" when address_in = 16#164D# else
		x"9601" when address_in = 16#164E# else
		x"940E" when address_in = 16#164F# else
		x"158B" when address_in = 16#1650# else
		x"2388" when address_in = 16#1651# else
		x"F019" when address_in = 16#1652# else
		x"2D99" when address_in = 16#1653# else
		x"2D88" when address_in = 16#1654# else
		x"C002" when address_in = 16#1655# else
		x"E080" when address_in = 16#1656# else
		x"E090" when address_in = 16#1657# else
		x"9628" when address_in = 16#1658# else
		x"B60F" when address_in = 16#1659# else
		x"94F8" when address_in = 16#165A# else
		x"BFDE" when address_in = 16#165B# else
		x"BE0F" when address_in = 16#165C# else
		x"BFCD" when address_in = 16#165D# else
		x"91DF" when address_in = 16#165E# else
		x"91CF" when address_in = 16#165F# else
		x"911F" when address_in = 16#1660# else
		x"910F" when address_in = 16#1661# else
		x"90FF" when address_in = 16#1662# else
		x"90EF" when address_in = 16#1663# else
		x"90DF" when address_in = 16#1664# else
		x"90CF" when address_in = 16#1665# else
		x"90BF" when address_in = 16#1666# else
		x"90AF" when address_in = 16#1667# else
		x"909F" when address_in = 16#1668# else
		x"908F" when address_in = 16#1669# else
		x"907F" when address_in = 16#166A# else
		x"9508" when address_in = 16#166B# else
		x"92CF" when address_in = 16#166C# else
		x"92DF" when address_in = 16#166D# else
		x"92EF" when address_in = 16#166E# else
		x"92FF" when address_in = 16#166F# else
		x"930F" when address_in = 16#1670# else
		x"931F" when address_in = 16#1671# else
		x"93CF" when address_in = 16#1672# else
		x"93DF" when address_in = 16#1673# else
		x"2EC6" when address_in = 16#1674# else
		x"2ED4" when address_in = 16#1675# else
		x"2FC2" when address_in = 16#1676# else
		x"940E" when address_in = 16#1677# else
		x"0B28" when address_in = 16#1678# else
		x"2FF9" when address_in = 16#1679# else
		x"2FE8" when address_in = 16#167A# else
		x"2B89" when address_in = 16#167B# else
		x"F429" when address_in = 16#167C# else
		x"940E" when address_in = 16#167D# else
		x"09DF" when address_in = 16#167E# else
		x"EE8A" when address_in = 16#167F# else
		x"EF9F" when address_in = 16#1680# else
		x"C039" when address_in = 16#1681# else
		x"8102" when address_in = 16#1682# else
		x"8113" when address_in = 16#1683# else
		x"80E6" when address_in = 16#1684# else
		x"80F7" when address_in = 16#1685# else
		x"2F2C" when address_in = 16#1686# else
		x"2D4D" when address_in = 16#1687# else
		x"2D6C" when address_in = 16#1688# else
		x"2F91" when address_in = 16#1689# else
		x"2F80" when address_in = 16#168A# else
		x"940E" when address_in = 16#168B# else
		x"15AB" when address_in = 16#168C# else
		x"27DD" when address_in = 16#168D# else
		x"9700" when address_in = 16#168E# else
		x"F039" when address_in = 16#168F# else
		x"0FCC" when address_in = 16#1690# else
		x"1FDD" when address_in = 16#1691# else
		x"0DCE" when address_in = 16#1692# else
		x"1DDF" when address_in = 16#1693# else
		x"8399" when address_in = 16#1694# else
		x"8388" when address_in = 16#1695# else
		x"C022" when address_in = 16#1696# else
		x"2FFD" when address_in = 16#1697# else
		x"2FEC" when address_in = 16#1698# else
		x"0FEC" when address_in = 16#1699# else
		x"1FFD" when address_in = 16#169A# else
		x"0DEE" when address_in = 16#169B# else
		x"1DFF" when address_in = 16#169C# else
		x"2F80" when address_in = 16#169D# else
		x"2F91" when address_in = 16#169E# else
		x"27AA" when address_in = 16#169F# else
		x"27BB" when address_in = 16#16A0# else
		x"0F88" when address_in = 16#16A1# else
		x"1F99" when address_in = 16#16A2# else
		x"1FAA" when address_in = 16#16A3# else
		x"1FBB" when address_in = 16#16A4# else
		x"E043" when address_in = 16#16A5# else
		x"0FCC" when address_in = 16#16A6# else
		x"1FDD" when address_in = 16#16A7# else
		x"954A" when address_in = 16#16A8# else
		x"F7E1" when address_in = 16#16A9# else
		x"962E" when address_in = 16#16AA# else
		x"2F2C" when address_in = 16#16AB# else
		x"2F3D" when address_in = 16#16AC# else
		x"2744" when address_in = 16#16AD# else
		x"2755" when address_in = 16#16AE# else
		x"0F82" when address_in = 16#16AF# else
		x"1F93" when address_in = 16#16B0# else
		x"1FA4" when address_in = 16#16B1# else
		x"1FB5" when address_in = 16#16B2# else
		x"95B6" when address_in = 16#16B3# else
		x"95A7" when address_in = 16#16B4# else
		x"9597" when address_in = 16#16B5# else
		x"9587" when address_in = 16#16B6# else
		x"8391" when address_in = 16#16B7# else
		x"8380" when address_in = 16#16B8# else
		x"E080" when address_in = 16#16B9# else
		x"E090" when address_in = 16#16BA# else
		x"91DF" when address_in = 16#16BB# else
		x"91CF" when address_in = 16#16BC# else
		x"911F" when address_in = 16#16BD# else
		x"910F" when address_in = 16#16BE# else
		x"90FF" when address_in = 16#16BF# else
		x"90EF" when address_in = 16#16C0# else
		x"90DF" when address_in = 16#16C1# else
		x"90CF" when address_in = 16#16C2# else
		x"9508" when address_in = 16#16C3# else
		x"930F" when address_in = 16#16C4# else
		x"931F" when address_in = 16#16C5# else
		x"2FB9" when address_in = 16#16C6# else
		x"2FA8" when address_in = 16#16C7# else
		x"2FF5" when address_in = 16#16C8# else
		x"2FE4" when address_in = 16#16C9# else
		x"2F86" when address_in = 16#16CA# else
		x"2799" when address_in = 16#16CB# else
		x"E073" when address_in = 16#16CC# else
		x"0F88" when address_in = 16#16CD# else
		x"1F99" when address_in = 16#16CE# else
		x"957A" when address_in = 16#16CF# else
		x"F7E1" when address_in = 16#16D0# else
		x"960E" when address_in = 16#16D1# else
		x"1780" when address_in = 16#16D2# else
		x"0791" when address_in = 16#16D3# else
		x"F170" when address_in = 16#16D4# else
		x"1501" when address_in = 16#16D5# else
		x"0511" when address_in = 16#16D6# else
		x"F449" when address_in = 16#16D7# else
		x"302E" when address_in = 16#16D8# else
		x"0531" when address_in = 16#16D9# else
		x"F030" when address_in = 16#16DA# else
		x"8584" when address_in = 16#16DB# else
		x"8595" when address_in = 16#16DC# else
		x"0F8A" when address_in = 16#16DD# else
		x"1F9B" when address_in = 16#16DE# else
		x"8795" when address_in = 16#16DF# else
		x"8784" when address_in = 16#16E0# else
		x"E070" when address_in = 16#16E1# else
		x"1776" when address_in = 16#16E2# else
		x"F4F8" when address_in = 16#16E3# else
		x"0F20" when address_in = 16#16E4# else
		x"1F31" when address_in = 16#16E5# else
		x"1BE0" when address_in = 16#16E6# else
		x"0BF1" when address_in = 16#16E7# else
		x"963E" when address_in = 16#16E8# else
		x"E040" when address_in = 16#16E9# else
		x"E050" when address_in = 16#16EA# else
		x"2F95" when address_in = 16#16EB# else
		x"2F84" when address_in = 16#16EC# else
		x"960E" when address_in = 16#16ED# else
		x"1780" when address_in = 16#16EE# else
		x"0791" when address_in = 16#16EF# else
		x"F060" when address_in = 16#16F0# else
		x"2F95" when address_in = 16#16F1# else
		x"2F84" when address_in = 16#16F2# else
		x"960F" when address_in = 16#16F3# else
		x"1782" when address_in = 16#16F4# else
		x"0793" when address_in = 16#16F5# else
		x"F430" when address_in = 16#16F6# else
		x"8180" when address_in = 16#16F7# else
		x"8191" when address_in = 16#16F8# else
		x"0F8A" when address_in = 16#16F9# else
		x"1F9B" when address_in = 16#16FA# else
		x"8391" when address_in = 16#16FB# else
		x"8380" when address_in = 16#16FC# else
		x"5F7F" when address_in = 16#16FD# else
		x"5F48" when address_in = 16#16FE# else
		x"4F5F" when address_in = 16#16FF# else
		x"9638" when address_in = 16#1700# else
		x"1776" when address_in = 16#1701# else
		x"F340" when address_in = 16#1702# else
		x"911F" when address_in = 16#1703# else
		x"910F" when address_in = 16#1704# else
		x"9508" when address_in = 16#1705# else
		x"930F" when address_in = 16#1706# else
		x"931F" when address_in = 16#1707# else
		x"2FB9" when address_in = 16#1708# else
		x"2FA8" when address_in = 16#1709# else
		x"2FF5" when address_in = 16#170A# else
		x"2FE4" when address_in = 16#170B# else
		x"2F86" when address_in = 16#170C# else
		x"2799" when address_in = 16#170D# else
		x"E043" when address_in = 16#170E# else
		x"0F88" when address_in = 16#170F# else
		x"1F99" when address_in = 16#1710# else
		x"954A" when address_in = 16#1711# else
		x"F7E1" when address_in = 16#1712# else
		x"960E" when address_in = 16#1713# else
		x"1780" when address_in = 16#1714# else
		x"0791" when address_in = 16#1715# else
		x"F170" when address_in = 16#1716# else
		x"1501" when address_in = 16#1717# else
		x"0511" when address_in = 16#1718# else
		x"F449" when address_in = 16#1719# else
		x"302E" when address_in = 16#171A# else
		x"0531" when address_in = 16#171B# else
		x"F030" when address_in = 16#171C# else
		x"8584" when address_in = 16#171D# else
		x"8595" when address_in = 16#171E# else
		x"1B8A" when address_in = 16#171F# else
		x"0B9B" when address_in = 16#1720# else
		x"8795" when address_in = 16#1721# else
		x"8784" when address_in = 16#1722# else
		x"E070" when address_in = 16#1723# else
		x"1776" when address_in = 16#1724# else
		x"F4F8" when address_in = 16#1725# else
		x"0F20" when address_in = 16#1726# else
		x"1F31" when address_in = 16#1727# else
		x"1BE0" when address_in = 16#1728# else
		x"0BF1" when address_in = 16#1729# else
		x"963E" when address_in = 16#172A# else
		x"E040" when address_in = 16#172B# else
		x"E050" when address_in = 16#172C# else
		x"2F95" when address_in = 16#172D# else
		x"2F84" when address_in = 16#172E# else
		x"960E" when address_in = 16#172F# else
		x"1780" when address_in = 16#1730# else
		x"0791" when address_in = 16#1731# else
		x"F060" when address_in = 16#1732# else
		x"2F95" when address_in = 16#1733# else
		x"2F84" when address_in = 16#1734# else
		x"960F" when address_in = 16#1735# else
		x"1782" when address_in = 16#1736# else
		x"0793" when address_in = 16#1737# else
		x"F430" when address_in = 16#1738# else
		x"8180" when address_in = 16#1739# else
		x"8191" when address_in = 16#173A# else
		x"1B8A" when address_in = 16#173B# else
		x"0B9B" when address_in = 16#173C# else
		x"8391" when address_in = 16#173D# else
		x"8380" when address_in = 16#173E# else
		x"5F7F" when address_in = 16#173F# else
		x"5F48" when address_in = 16#1740# else
		x"4F5F" when address_in = 16#1741# else
		x"9638" when address_in = 16#1742# else
		x"1776" when address_in = 16#1743# else
		x"F340" when address_in = 16#1744# else
		x"911F" when address_in = 16#1745# else
		x"910F" when address_in = 16#1746# else
		x"9508" when address_in = 16#1747# else
		x"925F" when address_in = 16#1748# else
		x"926F" when address_in = 16#1749# else
		x"927F" when address_in = 16#174A# else
		x"928F" when address_in = 16#174B# else
		x"929F" when address_in = 16#174C# else
		x"92AF" when address_in = 16#174D# else
		x"92BF" when address_in = 16#174E# else
		x"92CF" when address_in = 16#174F# else
		x"92DF" when address_in = 16#1750# else
		x"92EF" when address_in = 16#1751# else
		x"92FF" when address_in = 16#1752# else
		x"930F" when address_in = 16#1753# else
		x"931F" when address_in = 16#1754# else
		x"93CF" when address_in = 16#1755# else
		x"93DF" when address_in = 16#1756# else
		x"B7CD" when address_in = 16#1757# else
		x"B7DE" when address_in = 16#1758# else
		x"9724" when address_in = 16#1759# else
		x"B60F" when address_in = 16#175A# else
		x"94F8" when address_in = 16#175B# else
		x"BFDE" when address_in = 16#175C# else
		x"BE0F" when address_in = 16#175D# else
		x"BFCD" when address_in = 16#175E# else
		x"2EA8" when address_in = 16#175F# else
		x"2EB9" when address_in = 16#1760# else
		x"2FF9" when address_in = 16#1761# else
		x"2FE8" when address_in = 16#1762# else
		x"8126" when address_in = 16#1763# else
		x"8137" when address_in = 16#1764# else
		x"8182" when address_in = 16#1765# else
		x"8193" when address_in = 16#1766# else
		x"27AA" when address_in = 16#1767# else
		x"27BB" when address_in = 16#1768# else
		x"0F88" when address_in = 16#1769# else
		x"1F99" when address_in = 16#176A# else
		x"1FAA" when address_in = 16#176B# else
		x"1FBB" when address_in = 16#176C# else
		x"9603" when address_in = 16#176D# else
		x"1DA1" when address_in = 16#176E# else
		x"1DB1" when address_in = 16#176F# else
		x"BFAB" when address_in = 16#1770# else
		x"2FF9" when address_in = 16#1771# else
		x"2FE8" when address_in = 16#1772# else
		x"95D8" when address_in = 16#1773# else
		x"2C70" when address_in = 16#1774# else
		x"9601" when address_in = 16#1775# else
		x"1DA1" when address_in = 16#1776# else
		x"1DB1" when address_in = 16#1777# else
		x"BFAB" when address_in = 16#1778# else
		x"2FF9" when address_in = 16#1779# else
		x"2FE8" when address_in = 16#177A# else
		x"95D8" when address_in = 16#177B# else
		x"2C50" when address_in = 16#177C# else
		x"2466" when address_in = 16#177D# else
		x"1467" when address_in = 16#177E# else
		x"F008" when address_in = 16#177F# else
		x"C08E" when address_in = 16#1780# else
		x"E04E" when address_in = 16#1781# else
		x"E050" when address_in = 16#1782# else
		x"835A" when address_in = 16#1783# else
		x"8349" when address_in = 16#1784# else
		x"821C" when address_in = 16#1785# else
		x"821B" when address_in = 16#1786# else
		x"2EC2" when address_in = 16#1787# else
		x"2ED3" when address_in = 16#1788# else
		x"2DFB" when address_in = 16#1789# else
		x"2DEA" when address_in = 16#178A# else
		x"8082" when address_in = 16#178B# else
		x"8093" when address_in = 16#178C# else
		x"2CE8" when address_in = 16#178D# else
		x"2CF9" when address_in = 16#178E# else
		x"2700" when address_in = 16#178F# else
		x"2711" when address_in = 16#1790# else
		x"0CEE" when address_in = 16#1791# else
		x"1CFF" when address_in = 16#1792# else
		x"1F00" when address_in = 16#1793# else
		x"1F11" when address_in = 16#1794# else
		x"812B" when address_in = 16#1795# else
		x"813C" when address_in = 16#1796# else
		x"5E2C" when address_in = 16#1797# else
		x"4F3F" when address_in = 16#1798# else
		x"833C" when address_in = 16#1799# else
		x"832B" when address_in = 16#179A# else
		x"2F82" when address_in = 16#179B# else
		x"2F93" when address_in = 16#179C# else
		x"27AA" when address_in = 16#179D# else
		x"27BB" when address_in = 16#179E# else
		x"0D8E" when address_in = 16#179F# else
		x"1D9F" when address_in = 16#17A0# else
		x"1FA0" when address_in = 16#17A1# else
		x"1FB1" when address_in = 16#17A2# else
		x"BFAB" when address_in = 16#17A3# else
		x"2FF9" when address_in = 16#17A4# else
		x"2FE8" when address_in = 16#17A5# else
		x"95D8" when address_in = 16#17A6# else
		x"2D60" when address_in = 16#17A7# else
		x"5F2F" when address_in = 16#17A8# else
		x"4F3F" when address_in = 16#17A9# else
		x"2F82" when address_in = 16#17AA# else
		x"2F93" when address_in = 16#17AB# else
		x"27AA" when address_in = 16#17AC# else
		x"27BB" when address_in = 16#17AD# else
		x"5125" when address_in = 16#17AE# else
		x"4030" when address_in = 16#17AF# else
		x"833C" when address_in = 16#17B0# else
		x"832B" when address_in = 16#17B1# else
		x"0D8E" when address_in = 16#17B2# else
		x"1D9F" when address_in = 16#17B3# else
		x"1FA0" when address_in = 16#17B4# else
		x"1FB1" when address_in = 16#17B5# else
		x"BFAB" when address_in = 16#17B6# else
		x"2FF9" when address_in = 16#17B7# else
		x"2FE8" when address_in = 16#17B8# else
		x"95D8" when address_in = 16#17B9# else
		x"2D90" when address_in = 16#17BA# else
		x"2DFB" when address_in = 16#17BB# else
		x"2DEA" when address_in = 16#17BC# else
		x"8184" when address_in = 16#17BD# else
		x"1768" when address_in = 16#17BE# else
		x"F4A9" when address_in = 16#17BF# else
		x"E02E" when address_in = 16#17C0# else
		x"E030" when address_in = 16#17C1# else
		x"E040" when address_in = 16#17C2# else
		x"E050" when address_in = 16#17C3# else
		x"0EE2" when address_in = 16#17C4# else
		x"1EF3" when address_in = 16#17C5# else
		x"1F04" when address_in = 16#17C6# else
		x"1F15" when address_in = 16#17C7# else
		x"9516" when address_in = 16#17C8# else
		x"9507" when address_in = 16#17C9# else
		x"94F7" when address_in = 16#17CA# else
		x"94E7" when address_in = 16#17CB# else
		x"2D27" when address_in = 16#17CC# else
		x"0D25" when address_in = 16#17CD# else
		x"2D47" when address_in = 16#17CE# else
		x"2F69" when address_in = 16#17CF# else
		x"2D9F" when address_in = 16#17D0# else
		x"2D8E" when address_in = 16#17D1# else
		x"940E" when address_in = 16#17D2# else
		x"1544" when address_in = 16#17D3# else
		x"C008" when address_in = 16#17D4# else
		x"3F6F" when address_in = 16#17D5# else
		x"F041" when address_in = 16#17D6# else
		x"2D26" when address_in = 16#17D7# else
		x"2F49" when address_in = 16#17D8# else
		x"2D99" when address_in = 16#17D9# else
		x"2D88" when address_in = 16#17DA# else
		x"940E" when address_in = 16#17DB# else
		x"15AB" when address_in = 16#17DC# else
		x"9700" when address_in = 16#17DD# else
		x"F4C1" when address_in = 16#17DE# else
		x"2DFB" when address_in = 16#17DF# else
		x"2DEA" when address_in = 16#17E0# else
		x"8182" when address_in = 16#17E1# else
		x"8193" when address_in = 16#17E2# else
		x"27AA" when address_in = 16#17E3# else
		x"27BB" when address_in = 16#17E4# else
		x"0F88" when address_in = 16#17E5# else
		x"1F99" when address_in = 16#17E6# else
		x"1FAA" when address_in = 16#17E7# else
		x"1FBB" when address_in = 16#17E8# else
		x"8169" when address_in = 16#17E9# else
		x"817A" when address_in = 16#17EA# else
		x"2F26" when address_in = 16#17EB# else
		x"2F37" when address_in = 16#17EC# else
		x"2744" when address_in = 16#17ED# else
		x"2755" when address_in = 16#17EE# else
		x"0F82" when address_in = 16#17EF# else
		x"1F93" when address_in = 16#17F0# else
		x"1FA4" when address_in = 16#17F1# else
		x"1FB5" when address_in = 16#17F2# else
		x"95B6" when address_in = 16#17F3# else
		x"95A7" when address_in = 16#17F4# else
		x"9597" when address_in = 16#17F5# else
		x"9587" when address_in = 16#17F6# else
		x"2DFD" when address_in = 16#17F7# else
		x"2DEC" when address_in = 16#17F8# else
		x"8391" when address_in = 16#17F9# else
		x"8380" when address_in = 16#17FA# else
		x"9463" when address_in = 16#17FB# else
		x"E022" when address_in = 16#17FC# else
		x"E030" when address_in = 16#17FD# else
		x"0EC2" when address_in = 16#17FE# else
		x"1ED3" when address_in = 16#17FF# else
		x"814B" when address_in = 16#1800# else
		x"815C" when address_in = 16#1801# else
		x"5F48" when address_in = 16#1802# else
		x"4F5F" when address_in = 16#1803# else
		x"835C" when address_in = 16#1804# else
		x"834B" when address_in = 16#1805# else
		x"8169" when address_in = 16#1806# else
		x"817A" when address_in = 16#1807# else
		x"5F68" when address_in = 16#1808# else
		x"4F7F" when address_in = 16#1809# else
		x"837A" when address_in = 16#180A# else
		x"8369" when address_in = 16#180B# else
		x"1467" when address_in = 16#180C# else
		x"F408" when address_in = 16#180D# else
		x"CF7A" when address_in = 16#180E# else
		x"9624" when address_in = 16#180F# else
		x"B60F" when address_in = 16#1810# else
		x"94F8" when address_in = 16#1811# else
		x"BFDE" when address_in = 16#1812# else
		x"BE0F" when address_in = 16#1813# else
		x"BFCD" when address_in = 16#1814# else
		x"91DF" when address_in = 16#1815# else
		x"91CF" when address_in = 16#1816# else
		x"911F" when address_in = 16#1817# else
		x"910F" when address_in = 16#1818# else
		x"90FF" when address_in = 16#1819# else
		x"90EF" when address_in = 16#181A# else
		x"90DF" when address_in = 16#181B# else
		x"90CF" when address_in = 16#181C# else
		x"90BF" when address_in = 16#181D# else
		x"90AF" when address_in = 16#181E# else
		x"909F" when address_in = 16#181F# else
		x"908F" when address_in = 16#1820# else
		x"907F" when address_in = 16#1821# else
		x"906F" when address_in = 16#1822# else
		x"905F" when address_in = 16#1823# else
		x"9508" when address_in = 16#1824# else
		x"925F" when address_in = 16#1825# else
		x"926F" when address_in = 16#1826# else
		x"927F" when address_in = 16#1827# else
		x"928F" when address_in = 16#1828# else
		x"929F" when address_in = 16#1829# else
		x"92AF" when address_in = 16#182A# else
		x"92BF" when address_in = 16#182B# else
		x"92CF" when address_in = 16#182C# else
		x"92DF" when address_in = 16#182D# else
		x"92EF" when address_in = 16#182E# else
		x"92FF" when address_in = 16#182F# else
		x"930F" when address_in = 16#1830# else
		x"931F" when address_in = 16#1831# else
		x"93CF" when address_in = 16#1832# else
		x"93DF" when address_in = 16#1833# else
		x"B7CD" when address_in = 16#1834# else
		x"B7DE" when address_in = 16#1835# else
		x"976F" when address_in = 16#1836# else
		x"B60F" when address_in = 16#1837# else
		x"94F8" when address_in = 16#1838# else
		x"BFDE" when address_in = 16#1839# else
		x"BE0F" when address_in = 16#183A# else
		x"BFCD" when address_in = 16#183B# else
		x"879A" when address_in = 16#183C# else
		x"8789" when address_in = 16#183D# else
		x"876B" when address_in = 16#183E# else
		x"874C" when address_in = 16#183F# else
		x"872D" when address_in = 16#1840# else
		x"940E" when address_in = 16#1841# else
		x"0B61" when address_in = 16#1842# else
		x"879F" when address_in = 16#1843# else
		x"878E" when address_in = 16#1844# else
		x"8529" when address_in = 16#1845# else
		x"853A" when address_in = 16#1846# else
		x"2F82" when address_in = 16#1847# else
		x"2F93" when address_in = 16#1848# else
		x"27AA" when address_in = 16#1849# else
		x"27BB" when address_in = 16#184A# else
		x"0F88" when address_in = 16#184B# else
		x"1F99" when address_in = 16#184C# else
		x"1FAA" when address_in = 16#184D# else
		x"1FBB" when address_in = 16#184E# else
		x"854B" when address_in = 16#184F# else
		x"2F24" when address_in = 16#1850# else
		x"2733" when address_in = 16#1851# else
		x"E013" when address_in = 16#1852# else
		x"0F22" when address_in = 16#1853# else
		x"1F33" when address_in = 16#1854# else
		x"951A" when address_in = 16#1855# else
		x"F7E1" when address_in = 16#1856# else
		x"5F2A" when address_in = 16#1857# else
		x"4F3F" when address_in = 16#1858# else
		x"2744" when address_in = 16#1859# else
		x"2755" when address_in = 16#185A# else
		x"0F82" when address_in = 16#185B# else
		x"1F93" when address_in = 16#185C# else
		x"1FA4" when address_in = 16#185D# else
		x"1FB5" when address_in = 16#185E# else
		x"BFAB" when address_in = 16#185F# else
		x"2FF9" when address_in = 16#1860# else
		x"2FE8" when address_in = 16#1861# else
		x"95D8" when address_in = 16#1862# else
		x"2D60" when address_in = 16#1863# else
		x"8B69" when address_in = 16#1864# else
		x"8A18" when address_in = 16#1865# else
		x"8978" when address_in = 16#1866# else
		x"2FE7" when address_in = 16#1867# else
		x"27FF" when address_in = 16#1868# else
		x"0FEE" when address_in = 16#1869# else
		x"1FFF" when address_in = 16#186A# else
		x"858E" when address_in = 16#186B# else
		x"859F" when address_in = 16#186C# else
		x"0FE8" when address_in = 16#186D# else
		x"1FF9" when address_in = 16#186E# else
		x"80A0" when address_in = 16#186F# else
		x"80B1" when address_in = 16#1870# else
		x"14A1" when address_in = 16#1871# else
		x"04B1" when address_in = 16#1872# else
		x"F409" when address_in = 16#1873# else
		x"C17D" when address_in = 16#1874# else
		x"2DFB" when address_in = 16#1875# else
		x"2DEA" when address_in = 16#1876# else
		x"8182" when address_in = 16#1877# else
		x"8193" when address_in = 16#1878# else
		x"27AA" when address_in = 16#1879# else
		x"27BB" when address_in = 16#187A# else
		x"0F88" when address_in = 16#187B# else
		x"1F99" when address_in = 16#187C# else
		x"1FAA" when address_in = 16#187D# else
		x"1FBB" when address_in = 16#187E# else
		x"9603" when address_in = 16#187F# else
		x"1DA1" when address_in = 16#1880# else
		x"1DB1" when address_in = 16#1881# else
		x"BFAB" when address_in = 16#1882# else
		x"2FF9" when address_in = 16#1883# else
		x"2FE8" when address_in = 16#1884# else
		x"95D8" when address_in = 16#1885# else
		x"2D20" when address_in = 16#1886# else
		x"8B2A" when address_in = 16#1887# else
		x"8A1B" when address_in = 16#1888# else
		x"893B" when address_in = 16#1889# else
		x"1732" when address_in = 16#188A# else
		x"F008" when address_in = 16#188B# else
		x"C160" when address_in = 16#188C# else
		x"E06E" when address_in = 16#188D# else
		x"E070" when address_in = 16#188E# else
		x"8B7F" when address_in = 16#188F# else
		x"8B6E" when address_in = 16#1890# else
		x"8F79" when address_in = 16#1891# else
		x"8F68" when address_in = 16#1892# else
		x"8E1B" when address_in = 16#1893# else
		x"8E1A" when address_in = 16#1894# else
		x"E080" when address_in = 16#1895# else
		x"E090" when address_in = 16#1896# else
		x"8F9D" when address_in = 16#1897# else
		x"8F8C" when address_in = 16#1898# else
		x"8F9F" when address_in = 16#1899# else
		x"8F8E" when address_in = 16#189A# else
		x"2DFB" when address_in = 16#189B# else
		x"2DEA" when address_in = 16#189C# else
		x"8162" when address_in = 16#189D# else
		x"8173" when address_in = 16#189E# else
		x"2F26" when address_in = 16#189F# else
		x"2F37" when address_in = 16#18A0# else
		x"2744" when address_in = 16#18A1# else
		x"2755" when address_in = 16#18A2# else
		x"0F22" when address_in = 16#18A3# else
		x"1F33" when address_in = 16#18A4# else
		x"1F44" when address_in = 16#18A5# else
		x"1F55" when address_in = 16#18A6# else
		x"8D8A" when address_in = 16#18A7# else
		x"8D9B" when address_in = 16#18A8# else
		x"9644" when address_in = 16#18A9# else
		x"2FF9" when address_in = 16#18AA# else
		x"2FE8" when address_in = 16#18AB# else
		x"2F8E" when address_in = 16#18AC# else
		x"2F9F" when address_in = 16#18AD# else
		x"27AA" when address_in = 16#18AE# else
		x"27BB" when address_in = 16#18AF# else
		x"9774" when address_in = 16#18B0# else
		x"8FFB" when address_in = 16#18B1# else
		x"8FEA" when address_in = 16#18B2# else
		x"0F82" when address_in = 16#18B3# else
		x"1F93" when address_in = 16#18B4# else
		x"1FA4" when address_in = 16#18B5# else
		x"1FB5" when address_in = 16#18B6# else
		x"BFAB" when address_in = 16#18B7# else
		x"2FF9" when address_in = 16#18B8# else
		x"2FE8" when address_in = 16#18B9# else
		x"95D8" when address_in = 16#18BA# else
		x"2D80" when address_in = 16#18BB# else
		x"89F9" when address_in = 16#18BC# else
		x"178F" when address_in = 16#18BD# else
		x"F009" when address_in = 16#18BE# else
		x"C0E0" when address_in = 16#18BF# else
		x"8D6A" when address_in = 16#18C0# else
		x"8D7B" when address_in = 16#18C1# else
		x"5E6B" when address_in = 16#18C2# else
		x"4F7F" when address_in = 16#18C3# else
		x"2F86" when address_in = 16#18C4# else
		x"2F97" when address_in = 16#18C5# else
		x"27AA" when address_in = 16#18C6# else
		x"27BB" when address_in = 16#18C7# else
		x"5165" when address_in = 16#18C8# else
		x"4070" when address_in = 16#18C9# else
		x"8F7B" when address_in = 16#18CA# else
		x"8F6A" when address_in = 16#18CB# else
		x"0F28" when address_in = 16#18CC# else
		x"1F39" when address_in = 16#18CD# else
		x"1F4A" when address_in = 16#18CE# else
		x"1F5B" when address_in = 16#18CF# else
		x"BF4B" when address_in = 16#18D0# else
		x"2FF3" when address_in = 16#18D1# else
		x"2FE2" when address_in = 16#18D2# else
		x"95D8" when address_in = 16#18D3# else
		x"2D80" when address_in = 16#18D4# else
		x"852C" when address_in = 16#18D5# else
		x"854B" when address_in = 16#18D6# else
		x"2F68" when address_in = 16#18D7# else
		x"8589" when address_in = 16#18D8# else
		x"859A" when address_in = 16#18D9# else
		x"940E" when address_in = 16#18DA# else
		x"1544" when address_in = 16#18DB# else
		x"2E68" when address_in = 16#18DC# else
		x"2E79" when address_in = 16#18DD# else
		x"9700" when address_in = 16#18DE# else
		x"F409" when address_in = 16#18DF# else
		x"C0E9" when address_in = 16#18E0# else
		x"2DFB" when address_in = 16#18E1# else
		x"2DEA" when address_in = 16#18E2# else
		x"8006" when address_in = 16#18E3# else
		x"81F7" when address_in = 16#18E4# else
		x"2DE0" when address_in = 16#18E5# else
		x"8BFD" when address_in = 16#18E6# else
		x"8BEC" when address_in = 16#18E7# else
		x"2EE8" when address_in = 16#18E8# else
		x"2EF9" when address_in = 16#18E9# else
		x"2700" when address_in = 16#18EA# else
		x"2711" when address_in = 16#18EB# else
		x"0CEE" when address_in = 16#18EC# else
		x"1CFF" when address_in = 16#18ED# else
		x"1F00" when address_in = 16#18EE# else
		x"1F11" when address_in = 16#18EF# else
		x"2E8C" when address_in = 16#18F0# else
		x"2E9D" when address_in = 16#18F1# else
		x"9408" when address_in = 16#18F2# else
		x"1C81" when address_in = 16#18F3# else
		x"1C91" when address_in = 16#18F4# else
		x"8D6E" when address_in = 16#18F5# else
		x"8D7F" when address_in = 16#18F6# else
		x"5F60" when address_in = 16#18F7# else
		x"4F7F" when address_in = 16#18F8# else
		x"24CC" when address_in = 16#18F9# else
		x"24DD" when address_in = 16#18FA# else
		x"E053" when address_in = 16#18FB# else
		x"2E55" when address_in = 16#18FC# else
		x"2DFB" when address_in = 16#18FD# else
		x"2DEA" when address_in = 16#18FE# else
		x"8182" when address_in = 16#18FF# else
		x"8193" when address_in = 16#1900# else
		x"27AA" when address_in = 16#1901# else
		x"27BB" when address_in = 16#1902# else
		x"0F88" when address_in = 16#1903# else
		x"1F99" when address_in = 16#1904# else
		x"1FAA" when address_in = 16#1905# else
		x"1FBB" when address_in = 16#1906# else
		x"2F26" when address_in = 16#1907# else
		x"2F37" when address_in = 16#1908# else
		x"2744" when address_in = 16#1909# else
		x"2755" when address_in = 16#190A# else
		x"0F82" when address_in = 16#190B# else
		x"1F93" when address_in = 16#190C# else
		x"1FA4" when address_in = 16#190D# else
		x"1FB5" when address_in = 16#190E# else
		x"BFAB" when address_in = 16#190F# else
		x"2FF9" when address_in = 16#1910# else
		x"2FE8" when address_in = 16#1911# else
		x"95D8" when address_in = 16#1912# else
		x"2D80" when address_in = 16#1913# else
		x"2DB9" when address_in = 16#1914# else
		x"2DA8" when address_in = 16#1915# else
		x"938C" when address_in = 16#1916# else
		x"E0E2" when address_in = 16#1917# else
		x"E0F0" when address_in = 16#1918# else
		x"0ECE" when address_in = 16#1919# else
		x"1EDF" when address_in = 16#191A# else
		x"2D8C" when address_in = 16#191B# else
		x"2D9D" when address_in = 16#191C# else
		x"27AA" when address_in = 16#191D# else
		x"27BB" when address_in = 16#191E# else
		x"0D8E" when address_in = 16#191F# else
		x"1D9F" when address_in = 16#1920# else
		x"1FA0" when address_in = 16#1921# else
		x"1FB1" when address_in = 16#1922# else
		x"BFAB" when address_in = 16#1923# else
		x"2FF9" when address_in = 16#1924# else
		x"2FE8" when address_in = 16#1925# else
		x"95D8" when address_in = 16#1926# else
		x"2D80" when address_in = 16#1927# else
		x"2DF9" when address_in = 16#1928# else
		x"2DE8" when address_in = 16#1929# else
		x"8384" when address_in = 16#192A# else
		x"945A" when address_in = 16#192B# else
		x"9408" when address_in = 16#192C# else
		x"08C1" when address_in = 16#192D# else
		x"08D1" when address_in = 16#192E# else
		x"5F6F" when address_in = 16#192F# else
		x"4F7F" when address_in = 16#1930# else
		x"9408" when address_in = 16#1931# else
		x"1C81" when address_in = 16#1932# else
		x"1C91" when address_in = 16#1933# else
		x"FE57" when address_in = 16#1934# else
		x"CFC7" when address_in = 16#1935# else
		x"85FD" when address_in = 16#1936# else
		x"23FF" when address_in = 16#1937# else
		x"F0B9" when address_in = 16#1938# else
		x"2F6C" when address_in = 16#1939# else
		x"2F7D" when address_in = 16#193A# else
		x"5F6F" when address_in = 16#193B# else
		x"4F7F" when address_in = 16#193C# else
		x"2F8C" when address_in = 16#193D# else
		x"2F9D" when address_in = 16#193E# else
		x"9605" when address_in = 16#193F# else
		x"940E" when address_in = 16#1940# else
		x"158B" when address_in = 16#1941# else
		x"2388" when address_in = 16#1942# else
		x"F409" when address_in = 16#1943# else
		x"C085" when address_in = 16#1944# else
		x"8DEC" when address_in = 16#1945# else
		x"8DFD" when address_in = 16#1946# else
		x"0FEE" when address_in = 16#1947# else
		x"1FFF" when address_in = 16#1948# else
		x"892C" when address_in = 16#1949# else
		x"893D" when address_in = 16#194A# else
		x"0FE2" when address_in = 16#194B# else
		x"1FF3" when address_in = 16#194C# else
		x"8271" when address_in = 16#194D# else
		x"8260" when address_in = 16#194E# else
		x"C07A" when address_in = 16#194F# else
		x"8D0C" when address_in = 16#1950# else
		x"8D1D" when address_in = 16#1951# else
		x"0F00" when address_in = 16#1952# else
		x"1F11" when address_in = 16#1953# else
		x"896C" when address_in = 16#1954# else
		x"897D" when address_in = 16#1955# else
		x"0F06" when address_in = 16#1956# else
		x"1F17" when address_in = 16#1957# else
		x"2DFB" when address_in = 16#1958# else
		x"2DEA" when address_in = 16#1959# else
		x"8182" when address_in = 16#195A# else
		x"8193" when address_in = 16#195B# else
		x"27AA" when address_in = 16#195C# else
		x"27BB" when address_in = 16#195D# else
		x"0F88" when address_in = 16#195E# else
		x"1F99" when address_in = 16#195F# else
		x"1FAA" when address_in = 16#1960# else
		x"1FBB" when address_in = 16#1961# else
		x"8D68" when address_in = 16#1962# else
		x"8D79" when address_in = 16#1963# else
		x"2F26" when address_in = 16#1964# else
		x"2F37" when address_in = 16#1965# else
		x"2744" when address_in = 16#1966# else
		x"2755" when address_in = 16#1967# else
		x"0F82" when address_in = 16#1968# else
		x"1F93" when address_in = 16#1969# else
		x"1FA4" when address_in = 16#196A# else
		x"1FB5" when address_in = 16#196B# else
		x"95B6" when address_in = 16#196C# else
		x"95A7" when address_in = 16#196D# else
		x"9597" when address_in = 16#196E# else
		x"9587" when address_in = 16#196F# else
		x"2FF1" when address_in = 16#1970# else
		x"2FE0" when address_in = 16#1971# else
		x"8391" when address_in = 16#1972# else
		x"8380" when address_in = 16#1973# else
		x"C055" when address_in = 16#1974# else
		x"8DEC" when address_in = 16#1975# else
		x"8DFD" when address_in = 16#1976# else
		x"0FEE" when address_in = 16#1977# else
		x"1FFF" when address_in = 16#1978# else
		x"0FE4" when address_in = 16#1979# else
		x"1FF5" when address_in = 16#197A# else
		x"2F86" when address_in = 16#197B# else
		x"2F97" when address_in = 16#197C# else
		x"27AA" when address_in = 16#197D# else
		x"27BB" when address_in = 16#197E# else
		x"0F88" when address_in = 16#197F# else
		x"1F99" when address_in = 16#1980# else
		x"1FAA" when address_in = 16#1981# else
		x"1FBB" when address_in = 16#1982# else
		x"896E" when address_in = 16#1983# else
		x"897F" when address_in = 16#1984# else
		x"2F26" when address_in = 16#1985# else
		x"2F37" when address_in = 16#1986# else
		x"2744" when address_in = 16#1987# else
		x"2755" when address_in = 16#1988# else
		x"0F82" when address_in = 16#1989# else
		x"1F93" when address_in = 16#198A# else
		x"1FA4" when address_in = 16#198B# else
		x"1FB5" when address_in = 16#198C# else
		x"95B6" when address_in = 16#198D# else
		x"95A7" when address_in = 16#198E# else
		x"9597" when address_in = 16#198F# else
		x"9587" when address_in = 16#1990# else
		x"8391" when address_in = 16#1991# else
		x"8380" when address_in = 16#1992# else
		x"24EE" when address_in = 16#1993# else
		x"24FF" when address_in = 16#1994# else
		x"2D1F" when address_in = 16#1995# else
		x"2D0E" when address_in = 16#1996# else
		x"892B" when address_in = 16#1997# else
		x"E04A" when address_in = 16#1998# else
		x"E06C" when address_in = 16#1999# else
		x"2DFB" when address_in = 16#199A# else
		x"2DEA" when address_in = 16#199B# else
		x"8184" when address_in = 16#199C# else
		x"940E" when address_in = 16#199D# else
		x"0FD8" when address_in = 16#199E# else
		x"C02A" when address_in = 16#199F# else
		x"3F8F" when address_in = 16#19A0# else
		x"F541" when address_in = 16#19A1# else
		x"85FD" when address_in = 16#19A2# else
		x"23FF" when address_in = 16#19A3# else
		x"F529" when address_in = 16#19A4# else
		x"2DFB" when address_in = 16#19A5# else
		x"2DEA" when address_in = 16#19A6# else
		x"8146" when address_in = 16#19A7# else
		x"8157" when address_in = 16#19A8# else
		x"8DEC" when address_in = 16#19A9# else
		x"8DFD" when address_in = 16#19AA# else
		x"0FEE" when address_in = 16#19AB# else
		x"1FFF" when address_in = 16#19AC# else
		x"0FE4" when address_in = 16#19AD# else
		x"1FF5" when address_in = 16#19AE# else
		x"9001" when address_in = 16#19AF# else
		x"81F0" when address_in = 16#19B0# else
		x"2DE0" when address_in = 16#19B1# else
		x"852B" when address_in = 16#19B2# else
		x"853C" when address_in = 16#19B3# else
		x"1723" when address_in = 16#19B4# else
		x"F4A0" when address_in = 16#19B5# else
		x"2F82" when address_in = 16#19B6# else
		x"2799" when address_in = 16#19B7# else
		x"E0A3" when address_in = 16#19B8# else
		x"0F88" when address_in = 16#19B9# else
		x"1F99" when address_in = 16#19BA# else
		x"95AA" when address_in = 16#19BB# else
		x"F7E1" when address_in = 16#19BC# else
		x"85A9" when address_in = 16#19BD# else
		x"85BA" when address_in = 16#19BE# else
		x"0F8A" when address_in = 16#19BF# else
		x"1F9B" when address_in = 16#19C0# else
		x"178E" when address_in = 16#19C1# else
		x"079F" when address_in = 16#19C2# else
		x"F409" when address_in = 16#19C3# else
		x"CFB0" when address_in = 16#19C4# else
		x"5F2F" when address_in = 16#19C5# else
		x"9608" when address_in = 16#19C6# else
		x"85BC" when address_in = 16#19C7# else
		x"172B" when address_in = 16#19C8# else
		x"F3B8" when address_in = 16#19C9# else
		x"89EB" when address_in = 16#19CA# else
		x"5FEF" when address_in = 16#19CB# else
		x"8BEB" when address_in = 16#19CC# else
		x"8D2C" when address_in = 16#19CD# else
		x"8D3D" when address_in = 16#19CE# else
		x"5F2F" when address_in = 16#19CF# else
		x"4F3F" when address_in = 16#19D0# else
		x"8F3D" when address_in = 16#19D1# else
		x"8F2C" when address_in = 16#19D2# else
		x"8D6E" when address_in = 16#19D3# else
		x"8D7F" when address_in = 16#19D4# else
		x"5F68" when address_in = 16#19D5# else
		x"4F7F" when address_in = 16#19D6# else
		x"8F7F" when address_in = 16#19D7# else
		x"8F6E" when address_in = 16#19D8# else
		x"8D8A" when address_in = 16#19D9# else
		x"8D9B" when address_in = 16#19DA# else
		x"9608" when address_in = 16#19DB# else
		x"8F9B" when address_in = 16#19DC# else
		x"8F8A" when address_in = 16#19DD# else
		x"8DA8" when address_in = 16#19DE# else
		x"8DB9" when address_in = 16#19DF# else
		x"9618" when address_in = 16#19E0# else
		x"8FB9" when address_in = 16#19E1# else
		x"8FA8" when address_in = 16#19E2# else
		x"89EE" when address_in = 16#19E3# else
		x"89FF" when address_in = 16#19E4# else
		x"9638" when address_in = 16#19E5# else
		x"8BFF" when address_in = 16#19E6# else
		x"8BEE" when address_in = 16#19E7# else
		x"89FB" when address_in = 16#19E8# else
		x"892A" when address_in = 16#19E9# else
		x"17F2" when address_in = 16#19EA# else
		x"F408" when address_in = 16#19EB# else
		x"CEAE" when address_in = 16#19EC# else
		x"2DBB" when address_in = 16#19ED# else
		x"2DAA" when address_in = 16#19EE# else
		x"90AD" when address_in = 16#19EF# else
		x"90BC" when address_in = 16#19F0# else
		x"CE7F" when address_in = 16#19F1# else
		x"89B8" when address_in = 16#19F2# else
		x"5FBF" when address_in = 16#19F3# else
		x"8BB8" when address_in = 16#19F4# else
		x"30B4" when address_in = 16#19F5# else
		x"F408" when address_in = 16#19F6# else
		x"CE6E" when address_in = 16#19F7# else
		x"966F" when address_in = 16#19F8# else
		x"B60F" when address_in = 16#19F9# else
		x"94F8" when address_in = 16#19FA# else
		x"BFDE" when address_in = 16#19FB# else
		x"BE0F" when address_in = 16#19FC# else
		x"BFCD" when address_in = 16#19FD# else
		x"91DF" when address_in = 16#19FE# else
		x"91CF" when address_in = 16#19FF# else
		x"911F" when address_in = 16#1A00# else
		x"910F" when address_in = 16#1A01# else
		x"90FF" when address_in = 16#1A02# else
		x"90EF" when address_in = 16#1A03# else
		x"90DF" when address_in = 16#1A04# else
		x"90CF" when address_in = 16#1A05# else
		x"90BF" when address_in = 16#1A06# else
		x"90AF" when address_in = 16#1A07# else
		x"909F" when address_in = 16#1A08# else
		x"908F" when address_in = 16#1A09# else
		x"907F" when address_in = 16#1A0A# else
		x"906F" when address_in = 16#1A0B# else
		x"905F" when address_in = 16#1A0C# else
		x"9508" when address_in = 16#1A0D# else
		x"930F" when address_in = 16#1A0E# else
		x"931F" when address_in = 16#1A0F# else
		x"2F08" when address_in = 16#1A10# else
		x"2F19" when address_in = 16#1A11# else
		x"940E" when address_in = 16#1A12# else
		x"1748" when address_in = 16#1A13# else
		x"2FF1" when address_in = 16#1A14# else
		x"2FE0" when address_in = 16#1A15# else
		x"8182" when address_in = 16#1A16# else
		x"8193" when address_in = 16#1A17# else
		x"27AA" when address_in = 16#1A18# else
		x"27BB" when address_in = 16#1A19# else
		x"0F88" when address_in = 16#1A1A# else
		x"1F99" when address_in = 16#1A1B# else
		x"1FAA" when address_in = 16#1A1C# else
		x"1FBB" when address_in = 16#1A1D# else
		x"9604" when address_in = 16#1A1E# else
		x"1DA1" when address_in = 16#1A1F# else
		x"1DB1" when address_in = 16#1A20# else
		x"BFAB" when address_in = 16#1A21# else
		x"2FF9" when address_in = 16#1A22# else
		x"2FE8" when address_in = 16#1A23# else
		x"95D8" when address_in = 16#1A24# else
		x"2D40" when address_in = 16#1A25# else
		x"9701" when address_in = 16#1A26# else
		x"09A1" when address_in = 16#1A27# else
		x"09B1" when address_in = 16#1A28# else
		x"BFAB" when address_in = 16#1A29# else
		x"2FF9" when address_in = 16#1A2A# else
		x"2FE8" when address_in = 16#1A2B# else
		x"95D8" when address_in = 16#1A2C# else
		x"2D60" when address_in = 16#1A2D# else
		x"9703" when address_in = 16#1A2E# else
		x"09A1" when address_in = 16#1A2F# else
		x"09B1" when address_in = 16#1A30# else
		x"2344" when address_in = 16#1A31# else
		x"F059" when address_in = 16#1A32# else
		x"0F46" when address_in = 16#1A33# else
		x"960E" when address_in = 16#1A34# else
		x"1DA1" when address_in = 16#1A35# else
		x"1DB1" when address_in = 16#1A36# else
		x"95B6" when address_in = 16#1A37# else
		x"95A7" when address_in = 16#1A38# else
		x"9597" when address_in = 16#1A39# else
		x"9587" when address_in = 16#1A3A# else
		x"E021" when address_in = 16#1A3B# else
		x"940E" when address_in = 16#1A3C# else
		x"1825" when address_in = 16#1A3D# else
		x"E080" when address_in = 16#1A3E# else
		x"E090" when address_in = 16#1A3F# else
		x"911F" when address_in = 16#1A40# else
		x"910F" when address_in = 16#1A41# else
		x"9508" when address_in = 16#1A42# else
		x"92AF" when address_in = 16#1A43# else
		x"92BF" when address_in = 16#1A44# else
		x"92CF" when address_in = 16#1A45# else
		x"92DF" when address_in = 16#1A46# else
		x"92EF" when address_in = 16#1A47# else
		x"92FF" when address_in = 16#1A48# else
		x"930F" when address_in = 16#1A49# else
		x"931F" when address_in = 16#1A4A# else
		x"93CF" when address_in = 16#1A4B# else
		x"93DF" when address_in = 16#1A4C# else
		x"2FD9" when address_in = 16#1A4D# else
		x"2FC8" when address_in = 16#1A4E# else
		x"810E" when address_in = 16#1A4F# else
		x"811F" when address_in = 16#1A50# else
		x"818A" when address_in = 16#1A51# else
		x"819B" when address_in = 16#1A52# else
		x"27AA" when address_in = 16#1A53# else
		x"27BB" when address_in = 16#1A54# else
		x"0F88" when address_in = 16#1A55# else
		x"1F99" when address_in = 16#1A56# else
		x"1FAA" when address_in = 16#1A57# else
		x"1FBB" when address_in = 16#1A58# else
		x"9604" when address_in = 16#1A59# else
		x"1DA1" when address_in = 16#1A5A# else
		x"1DB1" when address_in = 16#1A5B# else
		x"BFAB" when address_in = 16#1A5C# else
		x"2FF9" when address_in = 16#1A5D# else
		x"2FE8" when address_in = 16#1A5E# else
		x"95D8" when address_in = 16#1A5F# else
		x"2D40" when address_in = 16#1A60# else
		x"9704" when address_in = 16#1A61# else
		x"09A1" when address_in = 16#1A62# else
		x"09B1" when address_in = 16#1A63# else
		x"2344" when address_in = 16#1A64# else
		x"F409" when address_in = 16#1A65# else
		x"C03D" when address_in = 16#1A66# else
		x"9603" when address_in = 16#1A67# else
		x"1DA1" when address_in = 16#1A68# else
		x"1DB1" when address_in = 16#1A69# else
		x"BFAB" when address_in = 16#1A6A# else
		x"2FF9" when address_in = 16#1A6B# else
		x"2FE8" when address_in = 16#1A6C# else
		x"95D8" when address_in = 16#1A6D# else
		x"2CD0" when address_in = 16#1A6E# else
		x"0D4D" when address_in = 16#1A6F# else
		x"960B" when address_in = 16#1A70# else
		x"1DA1" when address_in = 16#1A71# else
		x"1DB1" when address_in = 16#1A72# else
		x"95B6" when address_in = 16#1A73# else
		x"95A7" when address_in = 16#1A74# else
		x"9597" when address_in = 16#1A75# else
		x"9587" when address_in = 16#1A76# else
		x"E020" when address_in = 16#1A77# else
		x"2D6D" when address_in = 16#1A78# else
		x"940E" when address_in = 16#1A79# else
		x"1825" when address_in = 16#1A7A# else
		x"24CC" when address_in = 16#1A7B# else
		x"14CD" when address_in = 16#1A7C# else
		x"F530" when address_in = 16#1A7D# else
		x"2EA0" when address_in = 16#1A7E# else
		x"2EB1" when address_in = 16#1A7F# else
		x"2DFB" when address_in = 16#1A80# else
		x"2DEA" when address_in = 16#1A81# else
		x"9181" when address_in = 16#1A82# else
		x"9191" when address_in = 16#1A83# else
		x"2EAE" when address_in = 16#1A84# else
		x"2EBF" when address_in = 16#1A85# else
		x"27AA" when address_in = 16#1A86# else
		x"27BB" when address_in = 16#1A87# else
		x"0F88" when address_in = 16#1A88# else
		x"1F99" when address_in = 16#1A89# else
		x"1FAA" when address_in = 16#1A8A# else
		x"1FBB" when address_in = 16#1A8B# else
		x"9606" when address_in = 16#1A8C# else
		x"1DA1" when address_in = 16#1A8D# else
		x"1DB1" when address_in = 16#1A8E# else
		x"BFAB" when address_in = 16#1A8F# else
		x"2FF9" when address_in = 16#1A90# else
		x"2FE8" when address_in = 16#1A91# else
		x"95D8" when address_in = 16#1A92# else
		x"2D80" when address_in = 16#1A93# else
		x"812C" when address_in = 16#1A94# else
		x"1782" when address_in = 16#1A95# else
		x"F051" when address_in = 16#1A96# else
		x"3F8F" when address_in = 16#1A97# else
		x"F041" when address_in = 16#1A98# else
		x"24EE" when address_in = 16#1A99# else
		x"24FF" when address_in = 16#1A9A# else
		x"2D1F" when address_in = 16#1A9B# else
		x"2D0E" when address_in = 16#1A9C# else
		x"E04A" when address_in = 16#1A9D# else
		x"E06C" when address_in = 16#1A9E# else
		x"940E" when address_in = 16#1A9F# else
		x"0FD8" when address_in = 16#1AA0# else
		x"94C3" when address_in = 16#1AA1# else
		x"14CD" when address_in = 16#1AA2# else
		x"F2E0" when address_in = 16#1AA3# else
		x"E080" when address_in = 16#1AA4# else
		x"E090" when address_in = 16#1AA5# else
		x"91DF" when address_in = 16#1AA6# else
		x"91CF" when address_in = 16#1AA7# else
		x"911F" when address_in = 16#1AA8# else
		x"910F" when address_in = 16#1AA9# else
		x"90FF" when address_in = 16#1AAA# else
		x"90EF" when address_in = 16#1AAB# else
		x"90DF" when address_in = 16#1AAC# else
		x"90CF" when address_in = 16#1AAD# else
		x"90BF" when address_in = 16#1AAE# else
		x"90AF" when address_in = 16#1AAF# else
		x"9508" when address_in = 16#1AB0# else
		x"9508" when address_in = 16#1AB1# else
		x"EF8F" when address_in = 16#1AB2# else
		x"EF9F" when address_in = 16#1AB3# else
		x"9508" when address_in = 16#1AB4# else
		x"EF8F" when address_in = 16#1AB5# else
		x"EF9F" when address_in = 16#1AB6# else
		x"9508" when address_in = 16#1AB7# else
		x"EF6F" when address_in = 16#1AB8# else
		x"EF7F" when address_in = 16#1AB9# else
		x"EF8F" when address_in = 16#1ABA# else
		x"EF9F" when address_in = 16#1ABB# else
		x"9508" when address_in = 16#1ABC# else
		x"E080" when address_in = 16#1ABD# else
		x"E090" when address_in = 16#1ABE# else
		x"9508" when address_in = 16#1ABF# else
		x"930F" when address_in = 16#1AC0# else
		x"931F" when address_in = 16#1AC1# else
		x"93CF" when address_in = 16#1AC2# else
		x"93DF" when address_in = 16#1AC3# else
		x"2F08" when address_in = 16#1AC4# else
		x"2F19" when address_in = 16#1AC5# else
		x"2FD7" when address_in = 16#1AC6# else
		x"2FC6" when address_in = 16#1AC7# else
		x"2B67" when address_in = 16#1AC8# else
		x"F099" when address_in = 16#1AC9# else
		x"2F80" when address_in = 16#1ACA# else
		x"2F91" when address_in = 16#1ACB# else
		x"27AA" when address_in = 16#1ACC# else
		x"27BB" when address_in = 16#1ACD# else
		x"0F88" when address_in = 16#1ACE# else
		x"1F99" when address_in = 16#1ACF# else
		x"1FAA" when address_in = 16#1AD0# else
		x"1FBB" when address_in = 16#1AD1# else
		x"9606" when address_in = 16#1AD2# else
		x"1DA1" when address_in = 16#1AD3# else
		x"1DB1" when address_in = 16#1AD4# else
		x"BFAB" when address_in = 16#1AD5# else
		x"2FF9" when address_in = 16#1AD6# else
		x"2FE8" when address_in = 16#1AD7# else
		x"95D8" when address_in = 16#1AD8# else
		x"2D80" when address_in = 16#1AD9# else
		x"940E" when address_in = 16#1ADA# else
		x"0B54" when address_in = 16#1ADB# else
		x"8388" when address_in = 16#1ADC# else
		x"2F80" when address_in = 16#1ADD# else
		x"2F91" when address_in = 16#1ADE# else
		x"27AA" when address_in = 16#1ADF# else
		x"27BB" when address_in = 16#1AE0# else
		x"0F88" when address_in = 16#1AE1# else
		x"1F99" when address_in = 16#1AE2# else
		x"1FAA" when address_in = 16#1AE3# else
		x"1FBB" when address_in = 16#1AE4# else
		x"BFAB" when address_in = 16#1AE5# else
		x"2FF9" when address_in = 16#1AE6# else
		x"2FE8" when address_in = 16#1AE7# else
		x"95D8" when address_in = 16#1AE8# else
		x"2D80" when address_in = 16#1AE9# else
		x"B60B" when address_in = 16#1AEA# else
		x"9631" when address_in = 16#1AEB# else
		x"1C01" when address_in = 16#1AEC# else
		x"BE0B" when address_in = 16#1AED# else
		x"95D8" when address_in = 16#1AEE# else
		x"2D90" when address_in = 16#1AEF# else
		x"91DF" when address_in = 16#1AF0# else
		x"91CF" when address_in = 16#1AF1# else
		x"911F" when address_in = 16#1AF2# else
		x"910F" when address_in = 16#1AF3# else
		x"9508" when address_in = 16#1AF4# else
		x"92FF" when address_in = 16#1AF5# else
		x"930F" when address_in = 16#1AF6# else
		x"931F" when address_in = 16#1AF7# else
		x"2F08" when address_in = 16#1AF8# else
		x"2F19" when address_in = 16#1AF9# else
		x"B6FF" when address_in = 16#1AFA# else
		x"94F8" when address_in = 16#1AFB# else
		x"2F80" when address_in = 16#1AFC# else
		x"2F91" when address_in = 16#1AFD# else
		x"27AA" when address_in = 16#1AFE# else
		x"27BB" when address_in = 16#1AFF# else
		x"0F88" when address_in = 16#1B00# else
		x"1F99" when address_in = 16#1B01# else
		x"1FAA" when address_in = 16#1B02# else
		x"1FBB" when address_in = 16#1B03# else
		x"9606" when address_in = 16#1B04# else
		x"1DA1" when address_in = 16#1B05# else
		x"1DB1" when address_in = 16#1B06# else
		x"BFAB" when address_in = 16#1B07# else
		x"2FF9" when address_in = 16#1B08# else
		x"2FE8" when address_in = 16#1B09# else
		x"95D8" when address_in = 16#1B0A# else
		x"2D80" when address_in = 16#1B0B# else
		x"940E" when address_in = 16#1B0C# else
		x"0B54" when address_in = 16#1B0D# else
		x"91E0" when address_in = 16#1B0E# else
		x"0174" when address_in = 16#1B0F# else
		x"91F0" when address_in = 16#1B10# else
		x"0175" when address_in = 16#1B11# else
		x"8380" when address_in = 16#1B12# else
		x"9180" when address_in = 16#1B13# else
		x"0174" when address_in = 16#1B14# else
		x"9190" when address_in = 16#1B15# else
		x"0175" when address_in = 16#1B16# else
		x"9601" when address_in = 16#1B17# else
		x"9390" when address_in = 16#1B18# else
		x"0175" when address_in = 16#1B19# else
		x"9380" when address_in = 16#1B1A# else
		x"0174" when address_in = 16#1B1B# else
		x"BEFF" when address_in = 16#1B1C# else
		x"2F80" when address_in = 16#1B1D# else
		x"2F91" when address_in = 16#1B1E# else
		x"27AA" when address_in = 16#1B1F# else
		x"27BB" when address_in = 16#1B20# else
		x"0F88" when address_in = 16#1B21# else
		x"1F99" when address_in = 16#1B22# else
		x"1FAA" when address_in = 16#1B23# else
		x"1FBB" when address_in = 16#1B24# else
		x"BFAB" when address_in = 16#1B25# else
		x"2FF9" when address_in = 16#1B26# else
		x"2FE8" when address_in = 16#1B27# else
		x"95D8" when address_in = 16#1B28# else
		x"2D80" when address_in = 16#1B29# else
		x"B60B" when address_in = 16#1B2A# else
		x"9631" when address_in = 16#1B2B# else
		x"1C01" when address_in = 16#1B2C# else
		x"BE0B" when address_in = 16#1B2D# else
		x"95D8" when address_in = 16#1B2E# else
		x"2D90" when address_in = 16#1B2F# else
		x"911F" when address_in = 16#1B30# else
		x"910F" when address_in = 16#1B31# else
		x"90FF" when address_in = 16#1B32# else
		x"9508" when address_in = 16#1B33# else
		x"931F" when address_in = 16#1B34# else
		x"B71F" when address_in = 16#1B35# else
		x"94F8" when address_in = 16#1B36# else
		x"91E0" when address_in = 16#1B37# else
		x"0174" when address_in = 16#1B38# else
		x"91F0" when address_in = 16#1B39# else
		x"0175" when address_in = 16#1B3A# else
		x"9731" when address_in = 16#1B3B# else
		x"93F0" when address_in = 16#1B3C# else
		x"0175" when address_in = 16#1B3D# else
		x"93E0" when address_in = 16#1B3E# else
		x"0174" when address_in = 16#1B3F# else
		x"8180" when address_in = 16#1B40# else
		x"940E" when address_in = 16#1B41# else
		x"0B54" when address_in = 16#1B42# else
		x"BF1F" when address_in = 16#1B43# else
		x"911F" when address_in = 16#1B44# else
		x"9508" when address_in = 16#1B45# else
		x"92FF" when address_in = 16#1B46# else
		x"930F" when address_in = 16#1B47# else
		x"931F" when address_in = 16#1B48# else
		x"2EF8" when address_in = 16#1B49# else
		x"2F06" when address_in = 16#1B4A# else
		x"2F14" when address_in = 16#1B4B# else
		x"940E" when address_in = 16#1B4C# else
		x"0B5D" when address_in = 16#1B4D# else
		x"2F21" when address_in = 16#1B4E# else
		x"2F40" when address_in = 16#1B4F# else
		x"2D6F" when address_in = 16#1B50# else
		x"940E" when address_in = 16#1B51# else
		x"166C" when address_in = 16#1B52# else
		x"2799" when address_in = 16#1B53# else
		x"FD87" when address_in = 16#1B54# else
		x"9590" when address_in = 16#1B55# else
		x"911F" when address_in = 16#1B56# else
		x"910F" when address_in = 16#1B57# else
		x"90FF" when address_in = 16#1B58# else
		x"9508" when address_in = 16#1B59# else
		x"E087" when address_in = 16#1B5A# else
		x"E091" when address_in = 16#1B5B# else
		x"940E" when address_in = 16#1B5C# else
		x"2416" when address_in = 16#1B5D# else
		x"E08B" when address_in = 16#1B5E# else
		x"E091" when address_in = 16#1B5F# else
		x"940E" when address_in = 16#1B60# else
		x"2416" when address_in = 16#1B61# else
		x"E08F" when address_in = 16#1B62# else
		x"E091" when address_in = 16#1B63# else
		x"940E" when address_in = 16#1B64# else
		x"2416" when address_in = 16#1B65# else
		x"E183" when address_in = 16#1B66# else
		x"E091" when address_in = 16#1B67# else
		x"940E" when address_in = 16#1B68# else
		x"2416" when address_in = 16#1B69# else
		x"E080" when address_in = 16#1B6A# else
		x"E090" when address_in = 16#1B6B# else
		x"2F28" when address_in = 16#1B6C# else
		x"2F39" when address_in = 16#1B6D# else
		x"E043" when address_in = 16#1B6E# else
		x"2FF9" when address_in = 16#1B6F# else
		x"2FE8" when address_in = 16#1B70# else
		x"0FE2" when address_in = 16#1B71# else
		x"1FF3" when address_in = 16#1B72# else
		x"5EE9" when address_in = 16#1B73# else
		x"4FFE" when address_in = 16#1B74# else
		x"8215" when address_in = 16#1B75# else
		x"8214" when address_in = 16#1B76# else
		x"5041" when address_in = 16#1B77# else
		x"5F2F" when address_in = 16#1B78# else
		x"4F3F" when address_in = 16#1B79# else
		x"9605" when address_in = 16#1B7A# else
		x"FF47" when address_in = 16#1B7B# else
		x"CFF2" when address_in = 16#1B7C# else
		x"9508" when address_in = 16#1B7D# else
		x"93CF" when address_in = 16#1B7E# else
		x"93DF" when address_in = 16#1B7F# else
		x"2FD9" when address_in = 16#1B80# else
		x"2FC8" when address_in = 16#1B81# else
		x"81E8" when address_in = 16#1B82# else
		x"81F9" when address_in = 16#1B83# else
		x"9730" when address_in = 16#1B84# else
		x"F021" when address_in = 16#1B85# else
		x"818A" when address_in = 16#1B86# else
		x"819B" when address_in = 16#1B87# else
		x"2B89" when address_in = 16#1B88# else
		x"F419" when address_in = 16#1B89# else
		x"EE8A" when address_in = 16#1B8A# else
		x"EF9F" when address_in = 16#1B8B# else
		x"C01F" when address_in = 16#1B8C# else
		x"E081" when address_in = 16#1B8D# else
		x"30E7" when address_in = 16#1B8E# else
		x"07F8" when address_in = 16#1B8F# else
		x"F0A9" when address_in = 16#1B90# else
		x"852B" when address_in = 16#1B91# else
		x"853C" when address_in = 16#1B92# else
		x"854D" when address_in = 16#1B93# else
		x"855E" when address_in = 16#1B94# else
		x"1612" when address_in = 16#1B95# else
		x"0613" when address_in = 16#1B96# else
		x"0614" when address_in = 16#1B97# else
		x"0615" when address_in = 16#1B98# else
		x"F464" when address_in = 16#1B99# else
		x"8583" when address_in = 16#1B9A# else
		x"8594" when address_in = 16#1B9B# else
		x"85A5" when address_in = 16#1B9C# else
		x"85B6" when address_in = 16#1B9D# else
		x"0F82" when address_in = 16#1B9E# else
		x"1F93" when address_in = 16#1B9F# else
		x"1FA4" when address_in = 16#1BA0# else
		x"1FB5" when address_in = 16#1BA1# else
		x"8783" when address_in = 16#1BA2# else
		x"8794" when address_in = 16#1BA3# else
		x"87A5" when address_in = 16#1BA4# else
		x"87B6" when address_in = 16#1BA5# else
		x"2F8C" when address_in = 16#1BA6# else
		x"2F9D" when address_in = 16#1BA7# else
		x"940E" when address_in = 16#1BA8# else
		x"23D9" when address_in = 16#1BA9# else
		x"E080" when address_in = 16#1BAA# else
		x"E090" when address_in = 16#1BAB# else
		x"91DF" when address_in = 16#1BAC# else
		x"91CF" when address_in = 16#1BAD# else
		x"9508" when address_in = 16#1BAE# else
		x"92FF" when address_in = 16#1BAF# else
		x"930F" when address_in = 16#1BB0# else
		x"931F" when address_in = 16#1BB1# else
		x"93CF" when address_in = 16#1BB2# else
		x"93DF" when address_in = 16#1BB3# else
		x"2EF8" when address_in = 16#1BB4# else
		x"91C0" when address_in = 16#1BB5# else
		x"0107" when address_in = 16#1BB6# else
		x"91D0" when address_in = 16#1BB7# else
		x"0108" when address_in = 16#1BB8# else
		x"E081" when address_in = 16#1BB9# else
		x"30C7" when address_in = 16#1BBA# else
		x"07D8" when address_in = 16#1BBB# else
		x"F0E9" when address_in = 16#1BBC# else
		x"2F0C" when address_in = 16#1BBD# else
		x"2F1D" when address_in = 16#1BBE# else
		x"818D" when address_in = 16#1BBF# else
		x"158F" when address_in = 16#1BC0# else
		x"F4A1" when address_in = 16#1BC1# else
		x"800A" when address_in = 16#1BC2# else
		x"81DB" when address_in = 16#1BC3# else
		x"2DC0" when address_in = 16#1BC4# else
		x"2F91" when address_in = 16#1BC5# else
		x"2F80" when address_in = 16#1BC6# else
		x"940E" when address_in = 16#1BC7# else
		x"1B7E" when address_in = 16#1BC8# else
		x"B184" when address_in = 16#1BC9# else
		x"2799" when address_in = 16#1BCA# else
		x"718E" when address_in = 16#1BCB# else
		x"7090" when address_in = 16#1BCC# else
		x"9595" when address_in = 16#1BCD# else
		x"9587" when address_in = 16#1BCE# else
		x"9595" when address_in = 16#1BCF# else
		x"9587" when address_in = 16#1BD0# else
		x"2F68" when address_in = 16#1BD1# else
		x"2F91" when address_in = 16#1BD2# else
		x"2F80" when address_in = 16#1BD3# else
		x"940E" when address_in = 16#1BD4# else
		x"07EC" when address_in = 16#1BD5# else
		x"9009" when address_in = 16#1BD6# else
		x"81D8" when address_in = 16#1BD7# else
		x"2DC0" when address_in = 16#1BD8# else
		x"CFDF" when address_in = 16#1BD9# else
		x"91C0" when address_in = 16#1BDA# else
		x"010B" when address_in = 16#1BDB# else
		x"91D0" when address_in = 16#1BDC# else
		x"010C" when address_in = 16#1BDD# else
		x"E081" when address_in = 16#1BDE# else
		x"30CB" when address_in = 16#1BDF# else
		x"07D8" when address_in = 16#1BE0# else
		x"F0E9" when address_in = 16#1BE1# else
		x"2F0C" when address_in = 16#1BE2# else
		x"2F1D" when address_in = 16#1BE3# else
		x"818D" when address_in = 16#1BE4# else
		x"158F" when address_in = 16#1BE5# else
		x"F4A1" when address_in = 16#1BE6# else
		x"800A" when address_in = 16#1BE7# else
		x"81DB" when address_in = 16#1BE8# else
		x"2DC0" when address_in = 16#1BE9# else
		x"2F91" when address_in = 16#1BEA# else
		x"2F80" when address_in = 16#1BEB# else
		x"940E" when address_in = 16#1BEC# else
		x"23D9" when address_in = 16#1BED# else
		x"B184" when address_in = 16#1BEE# else
		x"2799" when address_in = 16#1BEF# else
		x"718E" when address_in = 16#1BF0# else
		x"7090" when address_in = 16#1BF1# else
		x"9595" when address_in = 16#1BF2# else
		x"9587" when address_in = 16#1BF3# else
		x"9595" when address_in = 16#1BF4# else
		x"9587" when address_in = 16#1BF5# else
		x"2F68" when address_in = 16#1BF6# else
		x"2F91" when address_in = 16#1BF7# else
		x"2F80" when address_in = 16#1BF8# else
		x"940E" when address_in = 16#1BF9# else
		x"07EC" when address_in = 16#1BFA# else
		x"9009" when address_in = 16#1BFB# else
		x"81D8" when address_in = 16#1BFC# else
		x"2DC0" when address_in = 16#1BFD# else
		x"CFDF" when address_in = 16#1BFE# else
		x"91C0" when address_in = 16#1BFF# else
		x"010F" when address_in = 16#1C00# else
		x"91D0" when address_in = 16#1C01# else
		x"0110" when address_in = 16#1C02# else
		x"E081" when address_in = 16#1C03# else
		x"30CF" when address_in = 16#1C04# else
		x"07D8" when address_in = 16#1C05# else
		x"F0E9" when address_in = 16#1C06# else
		x"2F0C" when address_in = 16#1C07# else
		x"2F1D" when address_in = 16#1C08# else
		x"818D" when address_in = 16#1C09# else
		x"158F" when address_in = 16#1C0A# else
		x"F4A1" when address_in = 16#1C0B# else
		x"800A" when address_in = 16#1C0C# else
		x"81DB" when address_in = 16#1C0D# else
		x"2DC0" when address_in = 16#1C0E# else
		x"2F91" when address_in = 16#1C0F# else
		x"2F80" when address_in = 16#1C10# else
		x"940E" when address_in = 16#1C11# else
		x"23D9" when address_in = 16#1C12# else
		x"B184" when address_in = 16#1C13# else
		x"2799" when address_in = 16#1C14# else
		x"718E" when address_in = 16#1C15# else
		x"7090" when address_in = 16#1C16# else
		x"9595" when address_in = 16#1C17# else
		x"9587" when address_in = 16#1C18# else
		x"9595" when address_in = 16#1C19# else
		x"9587" when address_in = 16#1C1A# else
		x"2F68" when address_in = 16#1C1B# else
		x"2F91" when address_in = 16#1C1C# else
		x"2F80" when address_in = 16#1C1D# else
		x"940E" when address_in = 16#1C1E# else
		x"07EC" when address_in = 16#1C1F# else
		x"9009" when address_in = 16#1C20# else
		x"81D8" when address_in = 16#1C21# else
		x"2DC0" when address_in = 16#1C22# else
		x"CFDF" when address_in = 16#1C23# else
		x"91C0" when address_in = 16#1C24# else
		x"0113" when address_in = 16#1C25# else
		x"91D0" when address_in = 16#1C26# else
		x"0114" when address_in = 16#1C27# else
		x"E081" when address_in = 16#1C28# else
		x"31C3" when address_in = 16#1C29# else
		x"07D8" when address_in = 16#1C2A# else
		x"F0E9" when address_in = 16#1C2B# else
		x"2F0C" when address_in = 16#1C2C# else
		x"2F1D" when address_in = 16#1C2D# else
		x"818D" when address_in = 16#1C2E# else
		x"158F" when address_in = 16#1C2F# else
		x"F4A1" when address_in = 16#1C30# else
		x"800A" when address_in = 16#1C31# else
		x"81DB" when address_in = 16#1C32# else
		x"2DC0" when address_in = 16#1C33# else
		x"2F91" when address_in = 16#1C34# else
		x"2F80" when address_in = 16#1C35# else
		x"940E" when address_in = 16#1C36# else
		x"23D9" when address_in = 16#1C37# else
		x"B184" when address_in = 16#1C38# else
		x"2799" when address_in = 16#1C39# else
		x"718E" when address_in = 16#1C3A# else
		x"7090" when address_in = 16#1C3B# else
		x"9595" when address_in = 16#1C3C# else
		x"9587" when address_in = 16#1C3D# else
		x"9595" when address_in = 16#1C3E# else
		x"9587" when address_in = 16#1C3F# else
		x"2F68" when address_in = 16#1C40# else
		x"2F91" when address_in = 16#1C41# else
		x"2F80" when address_in = 16#1C42# else
		x"940E" when address_in = 16#1C43# else
		x"07EC" when address_in = 16#1C44# else
		x"9009" when address_in = 16#1C45# else
		x"81D8" when address_in = 16#1C46# else
		x"2DC0" when address_in = 16#1C47# else
		x"CFDF" when address_in = 16#1C48# else
		x"E080" when address_in = 16#1C49# else
		x"E090" when address_in = 16#1C4A# else
		x"91DF" when address_in = 16#1C4B# else
		x"91CF" when address_in = 16#1C4C# else
		x"911F" when address_in = 16#1C4D# else
		x"910F" when address_in = 16#1C4E# else
		x"90FF" when address_in = 16#1C4F# else
		x"9508" when address_in = 16#1C50# else
		x"92BF" when address_in = 16#1C51# else
		x"92CF" when address_in = 16#1C52# else
		x"92DF" when address_in = 16#1C53# else
		x"92EF" when address_in = 16#1C54# else
		x"92FF" when address_in = 16#1C55# else
		x"930F" when address_in = 16#1C56# else
		x"931F" when address_in = 16#1C57# else
		x"93CF" when address_in = 16#1C58# else
		x"93DF" when address_in = 16#1C59# else
		x"B7CD" when address_in = 16#1C5A# else
		x"B7DE" when address_in = 16#1C5B# else
		x"9764" when address_in = 16#1C5C# else
		x"B60F" when address_in = 16#1C5D# else
		x"94F8" when address_in = 16#1C5E# else
		x"BFDE" when address_in = 16#1C5F# else
		x"BE0F" when address_in = 16#1C60# else
		x"BFCD" when address_in = 16#1C61# else
		x"2EB8" when address_in = 16#1C62# else
		x"2EE6" when address_in = 16#1C63# else
		x"E08A" when address_in = 16#1C64# else
		x"1786" when address_in = 16#1C65# else
		x"F418" when address_in = 16#1C66# else
		x"EE8A" when address_in = 16#1C67# else
		x"EF9F" when address_in = 16#1C68# else
		x"C053" when address_in = 16#1C69# else
		x"24FF" when address_in = 16#1C6A# else
		x"14FE" when address_in = 16#1C6B# else
		x"F5A0" when address_in = 16#1C6C# else
		x"2D0F" when address_in = 16#1C6D# else
		x"2711" when address_in = 16#1C6E# else
		x"0F00" when address_in = 16#1C6F# else
		x"1F11" when address_in = 16#1C70# else
		x"2ECC" when address_in = 16#1C71# else
		x"2EDD" when address_in = 16#1C72# else
		x"9408" when address_in = 16#1C73# else
		x"1CC1" when address_in = 16#1C74# else
		x"1CD1" when address_in = 16#1C75# else
		x"0D0C" when address_in = 16#1C76# else
		x"1D1D" when address_in = 16#1C77# else
		x"E064" when address_in = 16#1C78# else
		x"E180" when address_in = 16#1C79# else
		x"E090" when address_in = 16#1C7A# else
		x"940E" when address_in = 16#1C7B# else
		x"0640" when address_in = 16#1C7C# else
		x"2FF1" when address_in = 16#1C7D# else
		x"2FE0" when address_in = 16#1C7E# else
		x"8391" when address_in = 16#1C7F# else
		x"8380" when address_in = 16#1C80# else
		x"2B89" when address_in = 16#1C81# else
		x"F4E1" when address_in = 16#1C82# else
		x"24EE" when address_in = 16#1C83# else
		x"14EF" when address_in = 16#1C84# else
		x"F4B0" when address_in = 16#1C85# else
		x"2D1D" when address_in = 16#1C86# else
		x"2D0C" when address_in = 16#1C87# else
		x"B184" when address_in = 16#1C88# else
		x"2799" when address_in = 16#1C89# else
		x"718E" when address_in = 16#1C8A# else
		x"7090" when address_in = 16#1C8B# else
		x"9595" when address_in = 16#1C8C# else
		x"9587" when address_in = 16#1C8D# else
		x"9595" when address_in = 16#1C8E# else
		x"9587" when address_in = 16#1C8F# else
		x"2F68" when address_in = 16#1C90# else
		x"2FF1" when address_in = 16#1C91# else
		x"2FE0" when address_in = 16#1C92# else
		x"9181" when address_in = 16#1C93# else
		x"9191" when address_in = 16#1C94# else
		x"2F0E" when address_in = 16#1C95# else
		x"2F1F" when address_in = 16#1C96# else
		x"940E" when address_in = 16#1C97# else
		x"07EC" when address_in = 16#1C98# else
		x"94E3" when address_in = 16#1C99# else
		x"14EF" when address_in = 16#1C9A# else
		x"F360" when address_in = 16#1C9B# else
		x"EF84" when address_in = 16#1C9C# else
		x"EF9F" when address_in = 16#1C9D# else
		x"C01E" when address_in = 16#1C9E# else
		x"94F3" when address_in = 16#1C9F# else
		x"CFCA" when address_in = 16#1CA0# else
		x"24FF" when address_in = 16#1CA1# else
		x"14FE" when address_in = 16#1CA2# else
		x"F4B8" when address_in = 16#1CA3# else
		x"E000" when address_in = 16#1CA4# else
		x"E010" when address_in = 16#1CA5# else
		x"2FFD" when address_in = 16#1CA6# else
		x"2FEC" when address_in = 16#1CA7# else
		x"0FE0" when address_in = 16#1CA8# else
		x"1FF1" when address_in = 16#1CA9# else
		x"8001" when address_in = 16#1CAA# else
		x"81F2" when address_in = 16#1CAB# else
		x"2DE0" when address_in = 16#1CAC# else
		x"82B5" when address_in = 16#1CAD# else
		x"E082" when address_in = 16#1CAE# else
		x"8787" when address_in = 16#1CAF# else
		x"2F6E" when address_in = 16#1CB0# else
		x"2F7F" when address_in = 16#1CB1# else
		x"E08F" when address_in = 16#1CB2# else
		x"E091" when address_in = 16#1CB3# else
		x"940E" when address_in = 16#1CB4# else
		x"23D6" when address_in = 16#1CB5# else
		x"94F3" when address_in = 16#1CB6# else
		x"5F0E" when address_in = 16#1CB7# else
		x"4F1F" when address_in = 16#1CB8# else
		x"14FE" when address_in = 16#1CB9# else
		x"F358" when address_in = 16#1CBA# else
		x"E080" when address_in = 16#1CBB# else
		x"E090" when address_in = 16#1CBC# else
		x"9664" when address_in = 16#1CBD# else
		x"B60F" when address_in = 16#1CBE# else
		x"94F8" when address_in = 16#1CBF# else
		x"BFDE" when address_in = 16#1CC0# else
		x"BE0F" when address_in = 16#1CC1# else
		x"BFCD" when address_in = 16#1CC2# else
		x"91DF" when address_in = 16#1CC3# else
		x"91CF" when address_in = 16#1CC4# else
		x"911F" when address_in = 16#1CC5# else
		x"910F" when address_in = 16#1CC6# else
		x"90FF" when address_in = 16#1CC7# else
		x"90EF" when address_in = 16#1CC8# else
		x"90DF" when address_in = 16#1CC9# else
		x"90CF" when address_in = 16#1CCA# else
		x"90BF" when address_in = 16#1CCB# else
		x"9508" when address_in = 16#1CCC# else
		x"3065" when address_in = 16#1CCD# else
		x"0571" when address_in = 16#1CCE# else
		x"0581" when address_in = 16#1CCF# else
		x"0591" when address_in = 16#1CD0# else
		x"F42C" when address_in = 16#1CD1# else
		x"E065" when address_in = 16#1CD2# else
		x"E070" when address_in = 16#1CD3# else
		x"E080" when address_in = 16#1CD4# else
		x"E090" when address_in = 16#1CD5# else
		x"C009" when address_in = 16#1CD6# else
		x"3F6B" when address_in = 16#1CD7# else
		x"0571" when address_in = 16#1CD8# else
		x"0581" when address_in = 16#1CD9# else
		x"0591" when address_in = 16#1CDA# else
		x"F03C" when address_in = 16#1CDB# else
		x"EF6A" when address_in = 16#1CDC# else
		x"E070" when address_in = 16#1CDD# else
		x"E080" when address_in = 16#1CDE# else
		x"E090" when address_in = 16#1CDF# else
		x"940E" when address_in = 16#1CE0# else
		x"2D76" when address_in = 16#1CE1# else
		x"9508" when address_in = 16#1CE2# else
		x"2F86" when address_in = 16#1CE3# else
		x"2799" when address_in = 16#1CE4# else
		x"27AA" when address_in = 16#1CE5# else
		x"27BB" when address_in = 16#1CE6# else
		x"2F68" when address_in = 16#1CE7# else
		x"2F79" when address_in = 16#1CE8# else
		x"2F8A" when address_in = 16#1CE9# else
		x"2F9B" when address_in = 16#1CEA# else
		x"CFF4" when address_in = 16#1CEB# else
		x"927F" when address_in = 16#1CEC# else
		x"928F" when address_in = 16#1CED# else
		x"929F" when address_in = 16#1CEE# else
		x"92AF" when address_in = 16#1CEF# else
		x"92BF" when address_in = 16#1CF0# else
		x"92CF" when address_in = 16#1CF1# else
		x"92DF" when address_in = 16#1CF2# else
		x"92EF" when address_in = 16#1CF3# else
		x"92FF" when address_in = 16#1CF4# else
		x"930F" when address_in = 16#1CF5# else
		x"931F" when address_in = 16#1CF6# else
		x"93CF" when address_in = 16#1CF7# else
		x"93DF" when address_in = 16#1CF8# else
		x"B7CD" when address_in = 16#1CF9# else
		x"B7DE" when address_in = 16#1CFA# else
		x"972A" when address_in = 16#1CFB# else
		x"B60F" when address_in = 16#1CFC# else
		x"94F8" when address_in = 16#1CFD# else
		x"BFDE" when address_in = 16#1CFE# else
		x"BE0F" when address_in = 16#1CFF# else
		x"BFCD" when address_in = 16#1D00# else
		x"2E78" when address_in = 16#1D01# else
		x"EFFF" when address_in = 16#1D02# else
		x"2EAF" when address_in = 16#1D03# else
		x"2EBF" when address_in = 16#1D04# else
		x"2E8C" when address_in = 16#1D05# else
		x"2E9D" when address_in = 16#1D06# else
		x"9408" when address_in = 16#1D07# else
		x"1C81" when address_in = 16#1D08# else
		x"1C91" when address_in = 16#1D09# else
		x"90E0" when address_in = 16#1D0A# else
		x"0102" when address_in = 16#1D0B# else
		x"861A" when address_in = 16#1D0C# else
		x"8619" when address_in = 16#1D0D# else
		x"24CC" when address_in = 16#1D0E# else
		x"24DD" when address_in = 16#1D0F# else
		x"2D9D" when address_in = 16#1D10# else
		x"2D8C" when address_in = 16#1D11# else
		x"E0E3" when address_in = 16#1D12# else
		x"2EFE" when address_in = 16#1D13# else
		x"2D19" when address_in = 16#1D14# else
		x"2D08" when address_in = 16#1D15# else
		x"2FB1" when address_in = 16#1D16# else
		x"2FA0" when address_in = 16#1D17# else
		x"9611" when address_in = 16#1D18# else
		x"921C" when address_in = 16#1D19# else
		x"921E" when address_in = 16#1D1A# else
		x"2DFD" when address_in = 16#1D1B# else
		x"2DEC" when address_in = 16#1D1C# else
		x"0FE8" when address_in = 16#1D1D# else
		x"1FF9" when address_in = 16#1D1E# else
		x"5EE9" when address_in = 16#1D1F# else
		x"4FFE" when address_in = 16#1D20# else
		x"8144" when address_in = 16#1D21# else
		x"8155" when address_in = 16#1D22# else
		x"1541" when address_in = 16#1D23# else
		x"0551" when address_in = 16#1D24# else
		x"F149" when address_in = 16#1D25# else
		x"2D67" when address_in = 16#1D26# else
		x"2777" when address_in = 16#1D27# else
		x"8120" when address_in = 16#1D28# else
		x"8131" when address_in = 16#1D29# else
		x"1762" when address_in = 16#1D2A# else
		x"0773" when address_in = 16#1D2B# else
		x"F080" when address_in = 16#1D2C# else
		x"934D" when address_in = 16#1D2D# else
		x"935C" when address_in = 16#1D2E# else
		x"8142" when address_in = 16#1D2F# else
		x"8153" when address_in = 16#1D30# else
		x"1541" when address_in = 16#1D31# else
		x"0551" when address_in = 16#1D32# else
		x"F029" when address_in = 16#1D33# else
		x"1B46" when address_in = 16#1D34# else
		x"0B57" when address_in = 16#1D35# else
		x"0F24" when address_in = 16#1D36# else
		x"1F35" when address_in = 16#1D37# else
		x"C006" when address_in = 16#1D38# else
		x"8355" when address_in = 16#1D39# else
		x"8344" when address_in = 16#1D3A# else
		x"94EA" when address_in = 16#1D3B# else
		x"C012" when address_in = 16#1D3C# else
		x"1B26" when address_in = 16#1D3D# else
		x"0B37" when address_in = 16#1D3E# else
		x"8331" when address_in = 16#1D3F# else
		x"8320" when address_in = 16#1D40# else
		x"85E9" when address_in = 16#1D41# else
		x"85FA" when address_in = 16#1D42# else
		x"0FE8" when address_in = 16#1D43# else
		x"1FF9" when address_in = 16#1D44# else
		x"5EE9" when address_in = 16#1D45# else
		x"4FFE" when address_in = 16#1D46# else
		x"9001" when address_in = 16#1D47# else
		x"81F0" when address_in = 16#1D48# else
		x"2DE0" when address_in = 16#1D49# else
		x"15EA" when address_in = 16#1D4A# else
		x"05FB" when address_in = 16#1D4B# else
		x"F410" when address_in = 16#1D4C# else
		x"2EAE" when address_in = 16#1D4D# else
		x"2EBF" when address_in = 16#1D4E# else
		x"94FA" when address_in = 16#1D4F# else
		x"9601" when address_in = 16#1D50# else
		x"5F0E" when address_in = 16#1D51# else
		x"4F1F" when address_in = 16#1D52# else
		x"E0E5" when address_in = 16#1D53# else
		x"E0F0" when address_in = 16#1D54# else
		x"0ECE" when address_in = 16#1D55# else
		x"1EDF" when address_in = 16#1D56# else
		x"8529" when address_in = 16#1D57# else
		x"853A" when address_in = 16#1D58# else
		x"0F2E" when address_in = 16#1D59# else
		x"1F3F" when address_in = 16#1D5A# else
		x"873A" when address_in = 16#1D5B# else
		x"8729" when address_in = 16#1D5C# else
		x"FEF7" when address_in = 16#1D5D# else
		x"CFB7" when address_in = 16#1D5E# else
		x"92E0" when address_in = 16#1D5F# else
		x"0102" when address_in = 16#1D60# else
		x"E073" when address_in = 16#1D61# else
		x"2EF7" when address_in = 16#1D62# else
		x"2D19" when address_in = 16#1D63# else
		x"2D08" when address_in = 16#1D64# else
		x"2FB1" when address_in = 16#1D65# else
		x"2FA0" when address_in = 16#1D66# else
		x"91ED" when address_in = 16#1D67# else
		x"91FD" when address_in = 16#1D68# else
		x"2F0A" when address_in = 16#1D69# else
		x"2F1B" when address_in = 16#1D6A# else
		x"9730" when address_in = 16#1D6B# else
		x"F009" when address_in = 16#1D6C# else
		x"9509" when address_in = 16#1D6D# else
		x"94FA" when address_in = 16#1D6E# else
		x"FEF7" when address_in = 16#1D6F# else
		x"CFF4" when address_in = 16#1D70# else
		x"2D9B" when address_in = 16#1D71# else
		x"2D8A" when address_in = 16#1D72# else
		x"962A" when address_in = 16#1D73# else
		x"B60F" when address_in = 16#1D74# else
		x"94F8" when address_in = 16#1D75# else
		x"BFDE" when address_in = 16#1D76# else
		x"BE0F" when address_in = 16#1D77# else
		x"BFCD" when address_in = 16#1D78# else
		x"91DF" when address_in = 16#1D79# else
		x"91CF" when address_in = 16#1D7A# else
		x"911F" when address_in = 16#1D7B# else
		x"910F" when address_in = 16#1D7C# else
		x"90FF" when address_in = 16#1D7D# else
		x"90EF" when address_in = 16#1D7E# else
		x"90DF" when address_in = 16#1D7F# else
		x"90CF" when address_in = 16#1D80# else
		x"90BF" when address_in = 16#1D81# else
		x"90AF" when address_in = 16#1D82# else
		x"909F" when address_in = 16#1D83# else
		x"908F" when address_in = 16#1D84# else
		x"907F" when address_in = 16#1D85# else
		x"9508" when address_in = 16#1D86# else
		x"92EF" when address_in = 16#1D87# else
		x"92FF" when address_in = 16#1D88# else
		x"930F" when address_in = 16#1D89# else
		x"931F" when address_in = 16#1D8A# else
		x"93CF" when address_in = 16#1D8B# else
		x"2EE6" when address_in = 16#1D8C# else
		x"2EF7" when address_in = 16#1D8D# else
		x"2F08" when address_in = 16#1D8E# else
		x"2F19" when address_in = 16#1D8F# else
		x"B782" when address_in = 16#1D90# else
		x"2F28" when address_in = 16#1D91# else
		x"B7CF" when address_in = 16#1D92# else
		x"94F8" when address_in = 16#1D93# else
		x"2344" when address_in = 16#1D94# else
		x"F0A9" when address_in = 16#1D95# else
		x"9180" when address_in = 16#1D96# else
		x"0103" when address_in = 16#1D97# else
		x"9190" when address_in = 16#1D98# else
		x"0104" when address_in = 16#1D99# else
		x"91A0" when address_in = 16#1D9A# else
		x"0105" when address_in = 16#1D9B# else
		x"91B0" when address_in = 16#1D9C# else
		x"0106" when address_in = 16#1D9D# else
		x"0F82" when address_in = 16#1D9E# else
		x"1D91" when address_in = 16#1D9F# else
		x"1DA1" when address_in = 16#1DA0# else
		x"1DB1" when address_in = 16#1DA1# else
		x"9380" when address_in = 16#1DA2# else
		x"0103" when address_in = 16#1DA3# else
		x"9390" when address_in = 16#1DA4# else
		x"0104" when address_in = 16#1DA5# else
		x"93A0" when address_in = 16#1DA6# else
		x"0105" when address_in = 16#1DA7# else
		x"93B0" when address_in = 16#1DA8# else
		x"0106" when address_in = 16#1DA9# else
		x"C008" when address_in = 16#1DAA# else
		x"9210" when address_in = 16#1DAB# else
		x"0103" when address_in = 16#1DAC# else
		x"9210" when address_in = 16#1DAD# else
		x"0104" when address_in = 16#1DAE# else
		x"9210" when address_in = 16#1DAF# else
		x"0105" when address_in = 16#1DB0# else
		x"9210" when address_in = 16#1DB1# else
		x"0106" when address_in = 16#1DB2# else
		x"9180" when address_in = 16#1DB3# else
		x"0102" when address_in = 16#1DB4# else
		x"2388" when address_in = 16#1DB5# else
		x"F071" when address_in = 16#1DB6# else
		x"2F82" when address_in = 16#1DB7# else
		x"940E" when address_in = 16#1DB8# else
		x"1CEC" when address_in = 16#1DB9# else
		x"27AA" when address_in = 16#1DBA# else
		x"27BB" when address_in = 16#1DBB# else
		x"158E" when address_in = 16#1DBC# else
		x"059F" when address_in = 16#1DBD# else
		x"07A0" when address_in = 16#1DBE# else
		x"07B1" when address_in = 16#1DBF# else
		x"F424" when address_in = 16#1DC0# else
		x"2EE8" when address_in = 16#1DC1# else
		x"2EF9" when address_in = 16#1DC2# else
		x"2F0A" when address_in = 16#1DC3# else
		x"2F1B" when address_in = 16#1DC4# else
		x"2F91" when address_in = 16#1DC5# else
		x"2F80" when address_in = 16#1DC6# else
		x"2D7F" when address_in = 16#1DC7# else
		x"2D6E" when address_in = 16#1DC8# else
		x"940E" when address_in = 16#1DC9# else
		x"1CCD" when address_in = 16#1DCA# else
		x"BFCF" when address_in = 16#1DCB# else
		x"91CF" when address_in = 16#1DCC# else
		x"911F" when address_in = 16#1DCD# else
		x"910F" when address_in = 16#1DCE# else
		x"90FF" when address_in = 16#1DCF# else
		x"90EF" when address_in = 16#1DD0# else
		x"9508" when address_in = 16#1DD1# else
		x"92DF" when address_in = 16#1DD2# else
		x"92EF" when address_in = 16#1DD3# else
		x"92FF" when address_in = 16#1DD4# else
		x"930F" when address_in = 16#1DD5# else
		x"931F" when address_in = 16#1DD6# else
		x"93CF" when address_in = 16#1DD7# else
		x"93DF" when address_in = 16#1DD8# else
		x"2FD9" when address_in = 16#1DD9# else
		x"2FC8" when address_in = 16#1DDA# else
		x"2ED6" when address_in = 16#1DDB# else
		x"E087" when address_in = 16#1DDC# else
		x"E091" when address_in = 16#1DDD# else
		x"940E" when address_in = 16#1DDE# else
		x"241D" when address_in = 16#1DDF# else
		x"3081" when address_in = 16#1DE0# else
		x"F449" when address_in = 16#1DE1# else
		x"20DD" when address_in = 16#1DE2# else
		x"F409" when address_in = 16#1DE3# else
		x"C04E" when address_in = 16#1DE4# else
		x"E040" when address_in = 16#1DE5# else
		x"856B" when address_in = 16#1DE6# else
		x"857C" when address_in = 16#1DE7# else
		x"858D" when address_in = 16#1DE8# else
		x"859E" when address_in = 16#1DE9# else
		x"C046" when address_in = 16#1DEA# else
		x"B79F" when address_in = 16#1DEB# else
		x"94F8" when address_in = 16#1DEC# else
		x"B782" when address_in = 16#1DED# else
		x"90E0" when address_in = 16#1DEE# else
		x"0103" when address_in = 16#1DEF# else
		x"90F0" when address_in = 16#1DF0# else
		x"0104" when address_in = 16#1DF1# else
		x"9100" when address_in = 16#1DF2# else
		x"0105" when address_in = 16#1DF3# else
		x"9110" when address_in = 16#1DF4# else
		x"0106" when address_in = 16#1DF5# else
		x"0EE8" when address_in = 16#1DF6# else
		x"1CF1" when address_in = 16#1DF7# else
		x"1D01" when address_in = 16#1DF8# else
		x"1D11" when address_in = 16#1DF9# else
		x"BF9F" when address_in = 16#1DFA# else
		x"20DD" when address_in = 16#1DFB# else
		x"F061" when address_in = 16#1DFC# else
		x"858B" when address_in = 16#1DFD# else
		x"859C" when address_in = 16#1DFE# else
		x"85AD" when address_in = 16#1DFF# else
		x"85BE" when address_in = 16#1E00# else
		x"0D8E" when address_in = 16#1E01# else
		x"1D9F" when address_in = 16#1E02# else
		x"1FA0" when address_in = 16#1E03# else
		x"1FB1" when address_in = 16#1E04# else
		x"878B" when address_in = 16#1E05# else
		x"879C" when address_in = 16#1E06# else
		x"87AD" when address_in = 16#1E07# else
		x"87BE" when address_in = 16#1E08# else
		x"91E0" when address_in = 16#1E09# else
		x"0107" when address_in = 16#1E0A# else
		x"91F0" when address_in = 16#1E0B# else
		x"0108" when address_in = 16#1E0C# else
		x"852B" when address_in = 16#1E0D# else
		x"853C" when address_in = 16#1E0E# else
		x"854D" when address_in = 16#1E0F# else
		x"855E" when address_in = 16#1E10# else
		x"8583" when address_in = 16#1E11# else
		x"8594" when address_in = 16#1E12# else
		x"85A5" when address_in = 16#1E13# else
		x"85B6" when address_in = 16#1E14# else
		x"1728" when address_in = 16#1E15# else
		x"0739" when address_in = 16#1E16# else
		x"074A" when address_in = 16#1E17# else
		x"075B" when address_in = 16#1E18# else
		x"F57C" when address_in = 16#1E19# else
		x"1B82" when address_in = 16#1E1A# else
		x"0B93" when address_in = 16#1E1B# else
		x"0BA4" when address_in = 16#1E1C# else
		x"0BB5" when address_in = 16#1E1D# else
		x"8783" when address_in = 16#1E1E# else
		x"8794" when address_in = 16#1E1F# else
		x"87A5" when address_in = 16#1E20# else
		x"87B6" when address_in = 16#1E21# else
		x"20DD" when address_in = 16#1E22# else
		x"F079" when address_in = 16#1E23# else
		x"858B" when address_in = 16#1E24# else
		x"859C" when address_in = 16#1E25# else
		x"85AD" when address_in = 16#1E26# else
		x"85BE" when address_in = 16#1E27# else
		x"198E" when address_in = 16#1E28# else
		x"099F" when address_in = 16#1E29# else
		x"0BA0" when address_in = 16#1E2A# else
		x"0BB1" when address_in = 16#1E2B# else
		x"E041" when address_in = 16#1E2C# else
		x"2F68" when address_in = 16#1E2D# else
		x"2F79" when address_in = 16#1E2E# else
		x"2F8A" when address_in = 16#1E2F# else
		x"2F9B" when address_in = 16#1E30# else
		x"940E" when address_in = 16#1E31# else
		x"1D87" when address_in = 16#1E32# else
		x"2F6C" when address_in = 16#1E33# else
		x"2F7D" when address_in = 16#1E34# else
		x"E087" when address_in = 16#1E35# else
		x"E091" when address_in = 16#1E36# else
		x"940E" when address_in = 16#1E37# else
		x"23CF" when address_in = 16#1E38# else
		x"C032" when address_in = 16#1E39# else
		x"1B82" when address_in = 16#1E3A# else
		x"0B93" when address_in = 16#1E3B# else
		x"0BA4" when address_in = 16#1E3C# else
		x"0BB5" when address_in = 16#1E3D# else
		x"8783" when address_in = 16#1E3E# else
		x"8794" when address_in = 16#1E3F# else
		x"87A5" when address_in = 16#1E40# else
		x"87B6" when address_in = 16#1E41# else
		x"2F6C" when address_in = 16#1E42# else
		x"2F7D" when address_in = 16#1E43# else
		x"2F8E" when address_in = 16#1E44# else
		x"2F9F" when address_in = 16#1E45# else
		x"940E" when address_in = 16#1E46# else
		x"23B8" when address_in = 16#1E47# else
		x"C023" when address_in = 16#1E48# else
		x"E081" when address_in = 16#1E49# else
		x"30E7" when address_in = 16#1E4A# else
		x"07F8" when address_in = 16#1E4B# else
		x"F0C9" when address_in = 16#1E4C# else
		x"852B" when address_in = 16#1E4D# else
		x"853C" when address_in = 16#1E4E# else
		x"854D" when address_in = 16#1E4F# else
		x"855E" when address_in = 16#1E50# else
		x"8583" when address_in = 16#1E51# else
		x"8594" when address_in = 16#1E52# else
		x"85A5" when address_in = 16#1E53# else
		x"85B6" when address_in = 16#1E54# else
		x"1728" when address_in = 16#1E55# else
		x"0739" when address_in = 16#1E56# else
		x"074A" when address_in = 16#1E57# else
		x"075B" when address_in = 16#1E58# else
		x"F304" when address_in = 16#1E59# else
		x"1B28" when address_in = 16#1E5A# else
		x"0B39" when address_in = 16#1E5B# else
		x"0B4A" when address_in = 16#1E5C# else
		x"0B5B" when address_in = 16#1E5D# else
		x"872B" when address_in = 16#1E5E# else
		x"873C" when address_in = 16#1E5F# else
		x"874D" when address_in = 16#1E60# else
		x"875E" when address_in = 16#1E61# else
		x"9001" when address_in = 16#1E62# else
		x"81F0" when address_in = 16#1E63# else
		x"2DE0" when address_in = 16#1E64# else
		x"CFE3" when address_in = 16#1E65# else
		x"2F6C" when address_in = 16#1E66# else
		x"2F7D" when address_in = 16#1E67# else
		x"E087" when address_in = 16#1E68# else
		x"E091" when address_in = 16#1E69# else
		x"940E" when address_in = 16#1E6A# else
		x"23D6" when address_in = 16#1E6B# else
		x"91DF" when address_in = 16#1E6C# else
		x"91CF" when address_in = 16#1E6D# else
		x"911F" when address_in = 16#1E6E# else
		x"910F" when address_in = 16#1E6F# else
		x"90FF" when address_in = 16#1E70# else
		x"90EF" when address_in = 16#1E71# else
		x"90DF" when address_in = 16#1E72# else
		x"9508" when address_in = 16#1E73# else
		x"931F" when address_in = 16#1E74# else
		x"93CF" when address_in = 16#1E75# else
		x"2F18" when address_in = 16#1E76# else
		x"2FC6" when address_in = 16#1E77# else
		x"E087" when address_in = 16#1E78# else
		x"E091" when address_in = 16#1E79# else
		x"940E" when address_in = 16#1E7A# else
		x"241D" when address_in = 16#1E7B# else
		x"2388" when address_in = 16#1E7C# else
		x"F021" when address_in = 16#1E7D# else
		x"C014" when address_in = 16#1E7E# else
		x"2F8E" when address_in = 16#1E7F# else
		x"2F9F" when address_in = 16#1E80# else
		x"C013" when address_in = 16#1E81# else
		x"91E0" when address_in = 16#1E82# else
		x"0107" when address_in = 16#1E83# else
		x"91F0" when address_in = 16#1E84# else
		x"0108" when address_in = 16#1E85# else
		x"8185" when address_in = 16#1E86# else
		x"1781" when address_in = 16#1E87# else
		x"F419" when address_in = 16#1E88# else
		x"8186" when address_in = 16#1E89# else
		x"178C" when address_in = 16#1E8A# else
		x"F399" when address_in = 16#1E8B# else
		x"9001" when address_in = 16#1E8C# else
		x"81F0" when address_in = 16#1E8D# else
		x"2DE0" when address_in = 16#1E8E# else
		x"E081" when address_in = 16#1E8F# else
		x"30E7" when address_in = 16#1E90# else
		x"07F8" when address_in = 16#1E91# else
		x"F799" when address_in = 16#1E92# else
		x"E080" when address_in = 16#1E93# else
		x"E090" when address_in = 16#1E94# else
		x"91CF" when address_in = 16#1E95# else
		x"911F" when address_in = 16#1E96# else
		x"9508" when address_in = 16#1E97# else
		x"930F" when address_in = 16#1E98# else
		x"931F" when address_in = 16#1E99# else
		x"93CF" when address_in = 16#1E9A# else
		x"93DF" when address_in = 16#1E9B# else
		x"2F08" when address_in = 16#1E9C# else
		x"2F16" when address_in = 16#1E9D# else
		x"E183" when address_in = 16#1E9E# else
		x"E091" when address_in = 16#1E9F# else
		x"940E" when address_in = 16#1EA0# else
		x"241D" when address_in = 16#1EA1# else
		x"2388" when address_in = 16#1EA2# else
		x"F4C1" when address_in = 16#1EA3# else
		x"91C0" when address_in = 16#1EA4# else
		x"0113" when address_in = 16#1EA5# else
		x"91D0" when address_in = 16#1EA6# else
		x"0114" when address_in = 16#1EA7# else
		x"818D" when address_in = 16#1EA8# else
		x"1780" when address_in = 16#1EA9# else
		x"F451" when address_in = 16#1EAA# else
		x"818E" when address_in = 16#1EAB# else
		x"1781" when address_in = 16#1EAC# else
		x"F439" when address_in = 16#1EAD# else
		x"2F8C" when address_in = 16#1EAE# else
		x"2F9D" when address_in = 16#1EAF# else
		x"940E" when address_in = 16#1EB0# else
		x"23D9" when address_in = 16#1EB1# else
		x"2F8C" when address_in = 16#1EB2# else
		x"2F9D" when address_in = 16#1EB3# else
		x"C009" when address_in = 16#1EB4# else
		x"9009" when address_in = 16#1EB5# else
		x"81D8" when address_in = 16#1EB6# else
		x"2DC0" when address_in = 16#1EB7# else
		x"E081" when address_in = 16#1EB8# else
		x"31C3" when address_in = 16#1EB9# else
		x"07D8" when address_in = 16#1EBA# else
		x"F761" when address_in = 16#1EBB# else
		x"E080" when address_in = 16#1EBC# else
		x"E090" when address_in = 16#1EBD# else
		x"91DF" when address_in = 16#1EBE# else
		x"91CF" when address_in = 16#1EBF# else
		x"911F" when address_in = 16#1EC0# else
		x"910F" when address_in = 16#1EC1# else
		x"9508" when address_in = 16#1EC2# else
		x"930F" when address_in = 16#1EC3# else
		x"931F" when address_in = 16#1EC4# else
		x"93CF" when address_in = 16#1EC5# else
		x"93DF" when address_in = 16#1EC6# else
		x"2F08" when address_in = 16#1EC7# else
		x"2F16" when address_in = 16#1EC8# else
		x"E08B" when address_in = 16#1EC9# else
		x"E091" when address_in = 16#1ECA# else
		x"940E" when address_in = 16#1ECB# else
		x"241D" when address_in = 16#1ECC# else
		x"2388" when address_in = 16#1ECD# else
		x"F041" when address_in = 16#1ECE# else
		x"C018" when address_in = 16#1ECF# else
		x"2F8C" when address_in = 16#1ED0# else
		x"2F9D" when address_in = 16#1ED1# else
		x"940E" when address_in = 16#1ED2# else
		x"23D9" when address_in = 16#1ED3# else
		x"2F8C" when address_in = 16#1ED4# else
		x"2F9D" when address_in = 16#1ED5# else
		x"C013" when address_in = 16#1ED6# else
		x"91C0" when address_in = 16#1ED7# else
		x"010B" when address_in = 16#1ED8# else
		x"91D0" when address_in = 16#1ED9# else
		x"010C" when address_in = 16#1EDA# else
		x"818D" when address_in = 16#1EDB# else
		x"1780" when address_in = 16#1EDC# else
		x"F419" when address_in = 16#1EDD# else
		x"818E" when address_in = 16#1EDE# else
		x"1781" when address_in = 16#1EDF# else
		x"F379" when address_in = 16#1EE0# else
		x"9009" when address_in = 16#1EE1# else
		x"81D8" when address_in = 16#1EE2# else
		x"2DC0" when address_in = 16#1EE3# else
		x"E081" when address_in = 16#1EE4# else
		x"30CB" when address_in = 16#1EE5# else
		x"07D8" when address_in = 16#1EE6# else
		x"F799" when address_in = 16#1EE7# else
		x"E080" when address_in = 16#1EE8# else
		x"E090" when address_in = 16#1EE9# else
		x"91DF" when address_in = 16#1EEA# else
		x"91CF" when address_in = 16#1EEB# else
		x"911F" when address_in = 16#1EEC# else
		x"910F" when address_in = 16#1EED# else
		x"9508" when address_in = 16#1EEE# else
		x"930F" when address_in = 16#1EEF# else
		x"931F" when address_in = 16#1EF0# else
		x"93CF" when address_in = 16#1EF1# else
		x"93DF" when address_in = 16#1EF2# else
		x"2F08" when address_in = 16#1EF3# else
		x"2F16" when address_in = 16#1EF4# else
		x"940E" when address_in = 16#1EF5# else
		x"1E98" when address_in = 16#1EF6# else
		x"2FD9" when address_in = 16#1EF7# else
		x"2FC8" when address_in = 16#1EF8# else
		x"2B89" when address_in = 16#1EF9# else
		x"F469" when address_in = 16#1EFA# else
		x"2F61" when address_in = 16#1EFB# else
		x"2F80" when address_in = 16#1EFC# else
		x"940E" when address_in = 16#1EFD# else
		x"1E74" when address_in = 16#1EFE# else
		x"2FD9" when address_in = 16#1EFF# else
		x"2FC8" when address_in = 16#1F00# else
		x"9700" when address_in = 16#1F01# else
		x"F419" when address_in = 16#1F02# else
		x"EE8A" when address_in = 16#1F03# else
		x"EF9F" when address_in = 16#1F04# else
		x"C00A" when address_in = 16#1F05# else
		x"940E" when address_in = 16#1F06# else
		x"1B7E" when address_in = 16#1F07# else
		x"2F6C" when address_in = 16#1F08# else
		x"2F7D" when address_in = 16#1F09# else
		x"E08B" when address_in = 16#1F0A# else
		x"E091" when address_in = 16#1F0B# else
		x"940E" when address_in = 16#1F0C# else
		x"23D6" when address_in = 16#1F0D# else
		x"E080" when address_in = 16#1F0E# else
		x"E090" when address_in = 16#1F0F# else
		x"91DF" when address_in = 16#1F10# else
		x"91CF" when address_in = 16#1F11# else
		x"911F" when address_in = 16#1F12# else
		x"910F" when address_in = 16#1F13# else
		x"9508" when address_in = 16#1F14# else
		x"92FF" when address_in = 16#1F15# else
		x"930F" when address_in = 16#1F16# else
		x"931F" when address_in = 16#1F17# else
		x"93CF" when address_in = 16#1F18# else
		x"93DF" when address_in = 16#1F19# else
		x"2F18" when address_in = 16#1F1A# else
		x"2F06" when address_in = 16#1F1B# else
		x"2EF4" when address_in = 16#1F1C# else
		x"940E" when address_in = 16#1F1D# else
		x"1E98" when address_in = 16#1F1E# else
		x"2FD9" when address_in = 16#1F1F# else
		x"2FC8" when address_in = 16#1F20# else
		x"2B89" when address_in = 16#1F21# else
		x"F009" when address_in = 16#1F22# else
		x"C046" when address_in = 16#1F23# else
		x"2F60" when address_in = 16#1F24# else
		x"2F81" when address_in = 16#1F25# else
		x"940E" when address_in = 16#1F26# else
		x"1E74" when address_in = 16#1F27# else
		x"2FD9" when address_in = 16#1F28# else
		x"2FC8" when address_in = 16#1F29# else
		x"2B89" when address_in = 16#1F2A# else
		x"F031" when address_in = 16#1F2B# else
		x"2F60" when address_in = 16#1F2C# else
		x"2F81" when address_in = 16#1F2D# else
		x"940E" when address_in = 16#1F2E# else
		x"1EEF" when address_in = 16#1F2F# else
		x"82FC" when address_in = 16#1F30# else
		x"C03F" when address_in = 16#1F31# else
		x"2F60" when address_in = 16#1F32# else
		x"2F81" when address_in = 16#1F33# else
		x"940E" when address_in = 16#1F34# else
		x"1EC3" when address_in = 16#1F35# else
		x"2FD9" when address_in = 16#1F36# else
		x"2FC8" when address_in = 16#1F37# else
		x"2B89" when address_in = 16#1F38# else
		x"F571" when address_in = 16#1F39# else
		x"E08F" when address_in = 16#1F3A# else
		x"E091" when address_in = 16#1F3B# else
		x"940E" when address_in = 16#1F3C# else
		x"241D" when address_in = 16#1F3D# else
		x"2388" when address_in = 16#1F3E# else
		x"F041" when address_in = 16#1F3F# else
		x"C004" when address_in = 16#1F40# else
		x"2F8C" when address_in = 16#1F41# else
		x"2F9D" when address_in = 16#1F42# else
		x"940E" when address_in = 16#1F43# else
		x"23D9" when address_in = 16#1F44# else
		x"2F6C" when address_in = 16#1F45# else
		x"2F7D" when address_in = 16#1F46# else
		x"C010" when address_in = 16#1F47# else
		x"91C0" when address_in = 16#1F48# else
		x"010F" when address_in = 16#1F49# else
		x"91D0" when address_in = 16#1F4A# else
		x"0110" when address_in = 16#1F4B# else
		x"818D" when address_in = 16#1F4C# else
		x"1781" when address_in = 16#1F4D# else
		x"F391" when address_in = 16#1F4E# else
		x"9009" when address_in = 16#1F4F# else
		x"81D8" when address_in = 16#1F50# else
		x"2DC0" when address_in = 16#1F51# else
		x"E081" when address_in = 16#1F52# else
		x"30CF" when address_in = 16#1F53# else
		x"07D8" when address_in = 16#1F54# else
		x"F7B1" when address_in = 16#1F55# else
		x"E060" when address_in = 16#1F56# else
		x"E070" when address_in = 16#1F57# else
		x"2FD7" when address_in = 16#1F58# else
		x"2FC6" when address_in = 16#1F59# else
		x"2B67" when address_in = 16#1F5A# else
		x"F439" when address_in = 16#1F5B# else
		x"E064" when address_in = 16#1F5C# else
		x"E180" when address_in = 16#1F5D# else
		x"E090" when address_in = 16#1F5E# else
		x"940E" when address_in = 16#1F5F# else
		x"0640" when address_in = 16#1F60# else
		x"2FD9" when address_in = 16#1F61# else
		x"2FC8" when address_in = 16#1F62# else
		x"9720" when address_in = 16#1F63# else
		x"F419" when address_in = 16#1F64# else
		x"EF84" when address_in = 16#1F65# else
		x"EF9F" when address_in = 16#1F66# else
		x"C00B" when address_in = 16#1F67# else
		x"831D" when address_in = 16#1F68# else
		x"830E" when address_in = 16#1F69# else
		x"82FC" when address_in = 16#1F6A# else
		x"2F6C" when address_in = 16#1F6B# else
		x"2F7D" when address_in = 16#1F6C# else
		x"E08B" when address_in = 16#1F6D# else
		x"E091" when address_in = 16#1F6E# else
		x"940E" when address_in = 16#1F6F# else
		x"23D6" when address_in = 16#1F70# else
		x"E080" when address_in = 16#1F71# else
		x"E090" when address_in = 16#1F72# else
		x"91DF" when address_in = 16#1F73# else
		x"91CF" when address_in = 16#1F74# else
		x"911F" when address_in = 16#1F75# else
		x"910F" when address_in = 16#1F76# else
		x"90FF" when address_in = 16#1F77# else
		x"9508" when address_in = 16#1F78# else
		x"2FF9" when address_in = 16#1F79# else
		x"2FE8" when address_in = 16#1F7A# else
		x"8365" when address_in = 16#1F7B# else
		x"8346" when address_in = 16#1F7C# else
		x"8324" when address_in = 16#1F7D# else
		x"2F6E" when address_in = 16#1F7E# else
		x"2F7F" when address_in = 16#1F7F# else
		x"E08B" when address_in = 16#1F80# else
		x"E091" when address_in = 16#1F81# else
		x"940E" when address_in = 16#1F82# else
		x"23D6" when address_in = 16#1F83# else
		x"E080" when address_in = 16#1F84# else
		x"E090" when address_in = 16#1F85# else
		x"9508" when address_in = 16#1F86# else
		x"92EF" when address_in = 16#1F87# else
		x"92FF" when address_in = 16#1F88# else
		x"930F" when address_in = 16#1F89# else
		x"931F" when address_in = 16#1F8A# else
		x"2EE2" when address_in = 16#1F8B# else
		x"2EF3" when address_in = 16#1F8C# else
		x"2F04" when address_in = 16#1F8D# else
		x"2F15" when address_in = 16#1F8E# else
		x"940E" when address_in = 16#1F8F# else
		x"1EC3" when address_in = 16#1F90# else
		x"2FF9" when address_in = 16#1F91# else
		x"2FE8" when address_in = 16#1F92# else
		x"9700" when address_in = 16#1F93# else
		x"F419" when address_in = 16#1F94# else
		x"EE8A" when address_in = 16#1F95# else
		x"EF9F" when address_in = 16#1F96# else
		x"C00D" when address_in = 16#1F97# else
		x"82E7" when address_in = 16#1F98# else
		x"86F0" when address_in = 16#1F99# else
		x"8701" when address_in = 16#1F9A# else
		x"8712" when address_in = 16#1F9B# else
		x"86E3" when address_in = 16#1F9C# else
		x"86F4" when address_in = 16#1F9D# else
		x"8705" when address_in = 16#1F9E# else
		x"8716" when address_in = 16#1F9F# else
		x"E061" when address_in = 16#1FA0# else
		x"940E" when address_in = 16#1FA1# else
		x"1DD2" when address_in = 16#1FA2# else
		x"E080" when address_in = 16#1FA3# else
		x"E090" when address_in = 16#1FA4# else
		x"911F" when address_in = 16#1FA5# else
		x"910F" when address_in = 16#1FA6# else
		x"90FF" when address_in = 16#1FA7# else
		x"90EF" when address_in = 16#1FA8# else
		x"9508" when address_in = 16#1FA9# else
		x"930F" when address_in = 16#1FAA# else
		x"931F" when address_in = 16#1FAB# else
		x"2F08" when address_in = 16#1FAC# else
		x"2F16" when address_in = 16#1FAD# else
		x"940E" when address_in = 16#1FAE# else
		x"1EEF" when address_in = 16#1FAF# else
		x"2F61" when address_in = 16#1FB0# else
		x"2F80" when address_in = 16#1FB1# else
		x"940E" when address_in = 16#1FB2# else
		x"1EC3" when address_in = 16#1FB3# else
		x"2F28" when address_in = 16#1FB4# else
		x"2F39" when address_in = 16#1FB5# else
		x"2B89" when address_in = 16#1FB6# else
		x"F419" when address_in = 16#1FB7# else
		x"EE8A" when address_in = 16#1FB8# else
		x"EF9F" when address_in = 16#1FB9# else
		x"C00F" when address_in = 16#1FBA# else
		x"B184" when address_in = 16#1FBB# else
		x"2799" when address_in = 16#1FBC# else
		x"718E" when address_in = 16#1FBD# else
		x"7090" when address_in = 16#1FBE# else
		x"9595" when address_in = 16#1FBF# else
		x"9587" when address_in = 16#1FC0# else
		x"9595" when address_in = 16#1FC1# else
		x"9587" when address_in = 16#1FC2# else
		x"2F68" when address_in = 16#1FC3# else
		x"2F93" when address_in = 16#1FC4# else
		x"2F82" when address_in = 16#1FC5# else
		x"940E" when address_in = 16#1FC6# else
		x"07EC" when address_in = 16#1FC7# else
		x"E080" when address_in = 16#1FC8# else
		x"E090" when address_in = 16#1FC9# else
		x"911F" when address_in = 16#1FCA# else
		x"910F" when address_in = 16#1FCB# else
		x"9508" when address_in = 16#1FCC# else
		x"92CF" when address_in = 16#1FCD# else
		x"92DF" when address_in = 16#1FCE# else
		x"92EF" when address_in = 16#1FCF# else
		x"92FF" when address_in = 16#1FD0# else
		x"930F" when address_in = 16#1FD1# else
		x"931F" when address_in = 16#1FD2# else
		x"93CF" when address_in = 16#1FD3# else
		x"93DF" when address_in = 16#1FD4# else
		x"2EC8" when address_in = 16#1FD5# else
		x"2ED6" when address_in = 16#1FD6# else
		x"2EE2" when address_in = 16#1FD7# else
		x"2EF3" when address_in = 16#1FD8# else
		x"2F04" when address_in = 16#1FD9# else
		x"2F15" when address_in = 16#1FDA# else
		x"940E" when address_in = 16#1FDB# else
		x"1E98" when address_in = 16#1FDC# else
		x"2FD9" when address_in = 16#1FDD# else
		x"2FC8" when address_in = 16#1FDE# else
		x"2B89" when address_in = 16#1FDF# else
		x"F489" when address_in = 16#1FE0# else
		x"2D6D" when address_in = 16#1FE1# else
		x"2D8C" when address_in = 16#1FE2# else
		x"940E" when address_in = 16#1FE3# else
		x"1E74" when address_in = 16#1FE4# else
		x"2FD9" when address_in = 16#1FE5# else
		x"2FC8" when address_in = 16#1FE6# else
		x"9700" when address_in = 16#1FE7# else
		x"F019" when address_in = 16#1FE8# else
		x"940E" when address_in = 16#1FE9# else
		x"1B7E" when address_in = 16#1FEA# else
		x"C006" when address_in = 16#1FEB# else
		x"2D6D" when address_in = 16#1FEC# else
		x"2D8C" when address_in = 16#1FED# else
		x"940E" when address_in = 16#1FEE# else
		x"1EC3" when address_in = 16#1FEF# else
		x"2FD9" when address_in = 16#1FF0# else
		x"2FC8" when address_in = 16#1FF1# else
		x"9720" when address_in = 16#1FF2# else
		x"F419" when address_in = 16#1FF3# else
		x"EE8A" when address_in = 16#1FF4# else
		x"EF9F" when address_in = 16#1FF5# else
		x"C027" when address_in = 16#1FF6# else
		x"141E" when address_in = 16#1FF7# else
		x"041F" when address_in = 16#1FF8# else
		x"0610" when address_in = 16#1FF9# else
		x"0611" when address_in = 16#1FFA# else
		x"F024" when address_in = 16#1FFB# else
		x"80EF" when address_in = 16#1FFC# else
		x"84F8" when address_in = 16#1FFD# else
		x"8509" when address_in = 16#1FFE# else
		x"851A" when address_in = 16#1FFF# else
		x"E085" when address_in = 16#2000# else
		x"16E8" when address_in = 16#2001# else
		x"04F1" when address_in = 16#2002# else
		x"0501" when address_in = 16#2003# else
		x"0511" when address_in = 16#2004# else
		x"F44C" when address_in = 16#2005# else
		x"2F6C" when address_in = 16#2006# else
		x"2F7D" when address_in = 16#2007# else
		x"E08B" when address_in = 16#2008# else
		x"E091" when address_in = 16#2009# else
		x"940E" when address_in = 16#200A# else
		x"23D6" when address_in = 16#200B# else
		x"EF8F" when address_in = 16#200C# else
		x"EF9F" when address_in = 16#200D# else
		x"C00F" when address_in = 16#200E# else
		x"82EF" when address_in = 16#200F# else
		x"86F8" when address_in = 16#2010# else
		x"8709" when address_in = 16#2011# else
		x"871A" when address_in = 16#2012# else
		x"86EB" when address_in = 16#2013# else
		x"86FC" when address_in = 16#2014# else
		x"870D" when address_in = 16#2015# else
		x"871E" when address_in = 16#2016# else
		x"E061" when address_in = 16#2017# else
		x"2F8C" when address_in = 16#2018# else
		x"2F9D" when address_in = 16#2019# else
		x"940E" when address_in = 16#201A# else
		x"1DD2" when address_in = 16#201B# else
		x"E080" when address_in = 16#201C# else
		x"E090" when address_in = 16#201D# else
		x"91DF" when address_in = 16#201E# else
		x"91CF" when address_in = 16#201F# else
		x"911F" when address_in = 16#2020# else
		x"910F" when address_in = 16#2021# else
		x"90FF" when address_in = 16#2022# else
		x"90EF" when address_in = 16#2023# else
		x"90DF" when address_in = 16#2024# else
		x"90CF" when address_in = 16#2025# else
		x"9508" when address_in = 16#2026# else
		x"92CF" when address_in = 16#2027# else
		x"92DF" when address_in = 16#2028# else
		x"92EF" when address_in = 16#2029# else
		x"92FF" when address_in = 16#202A# else
		x"930F" when address_in = 16#202B# else
		x"931F" when address_in = 16#202C# else
		x"93CF" when address_in = 16#202D# else
		x"2F08" when address_in = 16#202E# else
		x"2EC4" when address_in = 16#202F# else
		x"2ED5" when address_in = 16#2030# else
		x"2EE6" when address_in = 16#2031# else
		x"2EF7" when address_in = 16#2032# else
		x"2F12" when address_in = 16#2033# else
		x"940E" when address_in = 16#2034# else
		x"0B5D" when address_in = 16#2035# else
		x"2FC8" when address_in = 16#2036# else
		x"2F41" when address_in = 16#2037# else
		x"2F60" when address_in = 16#2038# else
		x"940E" when address_in = 16#2039# else
		x"1F15" when address_in = 16#203A# else
		x"2388" when address_in = 16#203B# else
		x"F451" when address_in = 16#203C# else
		x"2D5F" when address_in = 16#203D# else
		x"2D4E" when address_in = 16#203E# else
		x"2D3D" when address_in = 16#203F# else
		x"2D2C" when address_in = 16#2040# else
		x"2F60" when address_in = 16#2041# else
		x"2F8C" when address_in = 16#2042# else
		x"940E" when address_in = 16#2043# else
		x"1F87" when address_in = 16#2044# else
		x"2388" when address_in = 16#2045# else
		x"F039" when address_in = 16#2046# else
		x"2F8C" when address_in = 16#2047# else
		x"940E" when address_in = 16#2048# else
		x"09FA" when address_in = 16#2049# else
		x"2799" when address_in = 16#204A# else
		x"FD87" when address_in = 16#204B# else
		x"9590" when address_in = 16#204C# else
		x"C002" when address_in = 16#204D# else
		x"E080" when address_in = 16#204E# else
		x"E090" when address_in = 16#204F# else
		x"91CF" when address_in = 16#2050# else
		x"911F" when address_in = 16#2051# else
		x"910F" when address_in = 16#2052# else
		x"90FF" when address_in = 16#2053# else
		x"90EF" when address_in = 16#2054# else
		x"90DF" when address_in = 16#2055# else
		x"90CF" when address_in = 16#2056# else
		x"9508" when address_in = 16#2057# else
		x"92DF" when address_in = 16#2058# else
		x"92EF" when address_in = 16#2059# else
		x"92FF" when address_in = 16#205A# else
		x"930F" when address_in = 16#205B# else
		x"931F" when address_in = 16#205C# else
		x"93CF" when address_in = 16#205D# else
		x"2ED8" when address_in = 16#205E# else
		x"2EE4" when address_in = 16#205F# else
		x"2EF5" when address_in = 16#2060# else
		x"2F06" when address_in = 16#2061# else
		x"2F17" when address_in = 16#2062# else
		x"940E" when address_in = 16#2063# else
		x"0B5D" when address_in = 16#2064# else
		x"2FC8" when address_in = 16#2065# else
		x"2F51" when address_in = 16#2066# else
		x"2F40" when address_in = 16#2067# else
		x"2D3F" when address_in = 16#2068# else
		x"2D2E" when address_in = 16#2069# else
		x"2D6D" when address_in = 16#206A# else
		x"940E" when address_in = 16#206B# else
		x"1FCD" when address_in = 16#206C# else
		x"2388" when address_in = 16#206D# else
		x"F039" when address_in = 16#206E# else
		x"2F8C" when address_in = 16#206F# else
		x"940E" when address_in = 16#2070# else
		x"09FA" when address_in = 16#2071# else
		x"2799" when address_in = 16#2072# else
		x"FD87" when address_in = 16#2073# else
		x"9590" when address_in = 16#2074# else
		x"C002" when address_in = 16#2075# else
		x"E080" when address_in = 16#2076# else
		x"E090" when address_in = 16#2077# else
		x"91CF" when address_in = 16#2078# else
		x"911F" when address_in = 16#2079# else
		x"910F" when address_in = 16#207A# else
		x"90FF" when address_in = 16#207B# else
		x"90EF" when address_in = 16#207C# else
		x"90DF" when address_in = 16#207D# else
		x"9508" when address_in = 16#207E# else
		x"931F" when address_in = 16#207F# else
		x"93CF" when address_in = 16#2080# else
		x"2F18" when address_in = 16#2081# else
		x"940E" when address_in = 16#2082# else
		x"0B5D" when address_in = 16#2083# else
		x"2FC8" when address_in = 16#2084# else
		x"2F61" when address_in = 16#2085# else
		x"940E" when address_in = 16#2086# else
		x"1EEF" when address_in = 16#2087# else
		x"2388" when address_in = 16#2088# else
		x"F431" when address_in = 16#2089# else
		x"2F61" when address_in = 16#208A# else
		x"2F8C" when address_in = 16#208B# else
		x"940E" when address_in = 16#208C# else
		x"1FAA" when address_in = 16#208D# else
		x"2388" when address_in = 16#208E# else
		x"F039" when address_in = 16#208F# else
		x"2F8C" when address_in = 16#2090# else
		x"940E" when address_in = 16#2091# else
		x"09FA" when address_in = 16#2092# else
		x"2799" when address_in = 16#2093# else
		x"FD87" when address_in = 16#2094# else
		x"9590" when address_in = 16#2095# else
		x"C002" when address_in = 16#2096# else
		x"E080" when address_in = 16#2097# else
		x"E090" when address_in = 16#2098# else
		x"91CF" when address_in = 16#2099# else
		x"911F" when address_in = 16#209A# else
		x"9508" when address_in = 16#209B# else
		x"92BF" when address_in = 16#209C# else
		x"92CF" when address_in = 16#209D# else
		x"92DF" when address_in = 16#209E# else
		x"92EF" when address_in = 16#209F# else
		x"92FF" when address_in = 16#20A0# else
		x"930F" when address_in = 16#20A1# else
		x"931F" when address_in = 16#20A2# else
		x"93CF" when address_in = 16#20A3# else
		x"93DF" when address_in = 16#20A4# else
		x"B78F" when address_in = 16#20A5# else
		x"94F8" when address_in = 16#20A6# else
		x"90E0" when address_in = 16#20A7# else
		x"0103" when address_in = 16#20A8# else
		x"90F0" when address_in = 16#20A9# else
		x"0104" when address_in = 16#20AA# else
		x"9100" when address_in = 16#20AB# else
		x"0105" when address_in = 16#20AC# else
		x"9110" when address_in = 16#20AD# else
		x"0106" when address_in = 16#20AE# else
		x"9210" when address_in = 16#20AF# else
		x"0103" when address_in = 16#20B0# else
		x"9210" when address_in = 16#20B1# else
		x"0104" when address_in = 16#20B2# else
		x"9210" when address_in = 16#20B3# else
		x"0105" when address_in = 16#20B4# else
		x"9210" when address_in = 16#20B5# else
		x"0106" when address_in = 16#20B6# else
		x"BF8F" when address_in = 16#20B7# else
		x"E087" when address_in = 16#20B8# else
		x"E091" when address_in = 16#20B9# else
		x"940E" when address_in = 16#20BA# else
		x"241D" when address_in = 16#20BB# else
		x"3081" when address_in = 16#20BC# else
		x"F409" when address_in = 16#20BD# else
		x"C07D" when address_in = 16#20BE# else
		x"91E0" when address_in = 16#20BF# else
		x"0107" when address_in = 16#20C0# else
		x"91F0" when address_in = 16#20C1# else
		x"0108" when address_in = 16#20C2# else
		x"E081" when address_in = 16#20C3# else
		x"30E7" when address_in = 16#20C4# else
		x"07F8" when address_in = 16#20C5# else
		x"F409" when address_in = 16#20C6# else
		x"C074" when address_in = 16#20C7# else
		x"8583" when address_in = 16#20C8# else
		x"8594" when address_in = 16#20C9# else
		x"85A5" when address_in = 16#20CA# else
		x"85B6" when address_in = 16#20CB# else
		x"2F28" when address_in = 16#20CC# else
		x"2F39" when address_in = 16#20CD# else
		x"2F4A" when address_in = 16#20CE# else
		x"2F5B" when address_in = 16#20CF# else
		x"192E" when address_in = 16#20D0# else
		x"093F" when address_in = 16#20D1# else
		x"0B40" when address_in = 16#20D2# else
		x"0B51" when address_in = 16#20D3# else
		x"158E" when address_in = 16#20D4# else
		x"059F" when address_in = 16#20D5# else
		x"07A0" when address_in = 16#20D6# else
		x"07B1" when address_in = 16#20D7# else
		x"F00C" when address_in = 16#20D8# else
		x"C0B7" when address_in = 16#20D9# else
		x"8723" when address_in = 16#20DA# else
		x"8734" when address_in = 16#20DB# else
		x"8745" when address_in = 16#20DC# else
		x"8756" when address_in = 16#20DD# else
		x"1AE8" when address_in = 16#20DE# else
		x"0AF9" when address_in = 16#20DF# else
		x"0B0A" when address_in = 16#20E0# else
		x"0B1B" when address_in = 16#20E1# else
		x"9001" when address_in = 16#20E2# else
		x"81F0" when address_in = 16#20E3# else
		x"2DE0" when address_in = 16#20E4# else
		x"CFDD" when address_in = 16#20E5# else
		x"91C0" when address_in = 16#20E6# else
		x"0107" when address_in = 16#20E7# else
		x"91D0" when address_in = 16#20E8# else
		x"0108" when address_in = 16#20E9# else
		x"858B" when address_in = 16#20EA# else
		x"859C" when address_in = 16#20EB# else
		x"85AD" when address_in = 16#20EC# else
		x"85BE" when address_in = 16#20ED# else
		x"1618" when address_in = 16#20EE# else
		x"0619" when address_in = 16#20EF# else
		x"061A" when address_in = 16#20F0# else
		x"061B" when address_in = 16#20F1# else
		x"F40C" when address_in = 16#20F2# else
		x"C05E" when address_in = 16#20F3# else
		x"80BD" when address_in = 16#20F4# else
		x"80CE" when address_in = 16#20F5# else
		x"E087" when address_in = 16#20F6# else
		x"E091" when address_in = 16#20F7# else
		x"940E" when address_in = 16#20F8# else
		x"2408" when address_in = 16#20F9# else
		x"818C" when address_in = 16#20FA# else
		x"FD81" when address_in = 16#20FB# else
		x"C003" when address_in = 16#20FC# else
		x"E4B0" when address_in = 16#20FD# else
		x"2EDB" when address_in = 16#20FE# else
		x"C001" when address_in = 16#20FF# else
		x"2ED1" when address_in = 16#2100# else
		x"FD80" when address_in = 16#2101# else
		x"C027" when address_in = 16#2102# else
		x"852B" when address_in = 16#2103# else
		x"853C" when address_in = 16#2104# else
		x"854D" when address_in = 16#2105# else
		x"855E" when address_in = 16#2106# else
		x"1612" when address_in = 16#2107# else
		x"0613" when address_in = 16#2108# else
		x"0614" when address_in = 16#2109# else
		x"0615" when address_in = 16#210A# else
		x"F0CC" when address_in = 16#210B# else
		x"80EF" when address_in = 16#210C# else
		x"84F8" when address_in = 16#210D# else
		x"8509" when address_in = 16#210E# else
		x"851A" when address_in = 16#210F# else
		x"2FB5" when address_in = 16#2110# else
		x"2FA4" when address_in = 16#2111# else
		x"2F93" when address_in = 16#2112# else
		x"2F82" when address_in = 16#2113# else
		x"0D8E" when address_in = 16#2114# else
		x"1D9F" when address_in = 16#2115# else
		x"1FA0" when address_in = 16#2116# else
		x"1FB1" when address_in = 16#2117# else
		x"2F28" when address_in = 16#2118# else
		x"2F39" when address_in = 16#2119# else
		x"2F4A" when address_in = 16#211A# else
		x"2F5B" when address_in = 16#211B# else
		x"1618" when address_in = 16#211C# else
		x"0619" when address_in = 16#211D# else
		x"061A" when address_in = 16#211E# else
		x"061B" when address_in = 16#211F# else
		x"F77C" when address_in = 16#2120# else
		x"878B" when address_in = 16#2121# else
		x"879C" when address_in = 16#2122# else
		x"87AD" when address_in = 16#2123# else
		x"87BE" when address_in = 16#2124# else
		x"2F6C" when address_in = 16#2125# else
		x"2F7D" when address_in = 16#2126# else
		x"E183" when address_in = 16#2127# else
		x"E091" when address_in = 16#2128# else
		x"C004" when address_in = 16#2129# else
		x"2F6C" when address_in = 16#212A# else
		x"2F7D" when address_in = 16#212B# else
		x"E08B" when address_in = 16#212C# else
		x"E091" when address_in = 16#212D# else
		x"940E" when address_in = 16#212E# else
		x"23D6" when address_in = 16#212F# else
		x"2D8D" when address_in = 16#2130# else
		x"2799" when address_in = 16#2131# else
		x"2EE8" when address_in = 16#2132# else
		x"2EF9" when address_in = 16#2133# else
		x"E000" when address_in = 16#2134# else
		x"E010" when address_in = 16#2135# else
		x"2D2C" when address_in = 16#2136# else
		x"E042" when address_in = 16#2137# else
		x"E064" when address_in = 16#2138# else
		x"2D8B" when address_in = 16#2139# else
		x"940E" when address_in = 16#213A# else
		x"0E67" when address_in = 16#213B# else
		x"E087" when address_in = 16#213C# else
		x"E091" when address_in = 16#213D# else
		x"940E" when address_in = 16#213E# else
		x"241D" when address_in = 16#213F# else
		x"2F18" when address_in = 16#2140# else
		x"2388" when address_in = 16#2141# else
		x"F409" when address_in = 16#2142# else
		x"CFA2" when address_in = 16#2143# else
		x"C00D" when address_in = 16#2144# else
		x"9100" when address_in = 16#2145# else
		x"0113" when address_in = 16#2146# else
		x"9110" when address_in = 16#2147# else
		x"0114" when address_in = 16#2148# else
		x"E183" when address_in = 16#2149# else
		x"E091" when address_in = 16#214A# else
		x"940E" when address_in = 16#214B# else
		x"2408" when address_in = 16#214C# else
		x"2F6C" when address_in = 16#214D# else
		x"2F91" when address_in = 16#214E# else
		x"2F80" when address_in = 16#214F# else
		x"940E" when address_in = 16#2150# else
		x"1DD2" when address_in = 16#2151# else
		x"E183" when address_in = 16#2152# else
		x"E091" when address_in = 16#2153# else
		x"940E" when address_in = 16#2154# else
		x"241D" when address_in = 16#2155# else
		x"2FC8" when address_in = 16#2156# else
		x"2388" when address_in = 16#2157# else
		x"F361" when address_in = 16#2158# else
		x"E087" when address_in = 16#2159# else
		x"E091" when address_in = 16#215A# else
		x"940E" when address_in = 16#215B# else
		x"241D" when address_in = 16#215C# else
		x"2388" when address_in = 16#215D# else
		x"F009" when address_in = 16#215E# else
		x"C03D" when address_in = 16#215F# else
		x"91E0" when address_in = 16#2160# else
		x"0107" when address_in = 16#2161# else
		x"91F0" when address_in = 16#2162# else
		x"0108" when address_in = 16#2163# else
		x"B7CF" when address_in = 16#2164# else
		x"94F8" when address_in = 16#2165# else
		x"B782" when address_in = 16#2166# else
		x"9120" when address_in = 16#2167# else
		x"0103" when address_in = 16#2168# else
		x"9130" when address_in = 16#2169# else
		x"0104" when address_in = 16#216A# else
		x"9140" when address_in = 16#216B# else
		x"0105" when address_in = 16#216C# else
		x"9150" when address_in = 16#216D# else
		x"0106" when address_in = 16#216E# else
		x"1B28" when address_in = 16#216F# else
		x"0931" when address_in = 16#2170# else
		x"0941" when address_in = 16#2171# else
		x"0951" when address_in = 16#2172# else
		x"84E3" when address_in = 16#2173# else
		x"84F4" when address_in = 16#2174# else
		x"8505" when address_in = 16#2175# else
		x"8516" when address_in = 16#2176# else
		x"2FB1" when address_in = 16#2177# else
		x"2FA0" when address_in = 16#2178# else
		x"2D9F" when address_in = 16#2179# else
		x"2D8E" when address_in = 16#217A# else
		x"1B82" when address_in = 16#217B# else
		x"0B93" when address_in = 16#217C# else
		x"0BA4" when address_in = 16#217D# else
		x"0BB5" when address_in = 16#217E# else
		x"1618" when address_in = 16#217F# else
		x"0619" when address_in = 16#2180# else
		x"061A" when address_in = 16#2181# else
		x"061B" when address_in = 16#2182# else
		x"F494" when address_in = 16#2183# else
		x"BFCF" when address_in = 16#2184# else
		x"1AE2" when address_in = 16#2185# else
		x"0AF3" when address_in = 16#2186# else
		x"0B04" when address_in = 16#2187# else
		x"0B15" when address_in = 16#2188# else
		x"E041" when address_in = 16#2189# else
		x"2F91" when address_in = 16#218A# else
		x"2F80" when address_in = 16#218B# else
		x"2D7F" when address_in = 16#218C# else
		x"2D6E" when address_in = 16#218D# else
		x"940E" when address_in = 16#218E# else
		x"1D87" when address_in = 16#218F# else
		x"C016" when address_in = 16#2190# else
		x"8723" when address_in = 16#2191# else
		x"8734" when address_in = 16#2192# else
		x"8745" when address_in = 16#2193# else
		x"8756" when address_in = 16#2194# else
		x"CFA6" when address_in = 16#2195# else
		x"BFCF" when address_in = 16#2196# else
		x"E96C" when address_in = 16#2197# else
		x"E270" when address_in = 16#2198# else
		x"E080" when address_in = 16#2199# else
		x"940E" when address_in = 16#219A# else
		x"0B1A" when address_in = 16#219B# else
		x"C00A" when address_in = 16#219C# else
		x"B7CF" when address_in = 16#219D# else
		x"94F8" when address_in = 16#219E# else
		x"E040" when address_in = 16#219F# else
		x"EF6A" when address_in = 16#21A0# else
		x"E070" when address_in = 16#21A1# else
		x"E080" when address_in = 16#21A2# else
		x"E090" when address_in = 16#21A3# else
		x"940E" when address_in = 16#21A4# else
		x"1D87" when address_in = 16#21A5# else
		x"BFCF" when address_in = 16#21A6# else
		x"91DF" when address_in = 16#21A7# else
		x"91CF" when address_in = 16#21A8# else
		x"911F" when address_in = 16#21A9# else
		x"910F" when address_in = 16#21AA# else
		x"90FF" when address_in = 16#21AB# else
		x"90EF" when address_in = 16#21AC# else
		x"90DF" when address_in = 16#21AD# else
		x"90CF" when address_in = 16#21AE# else
		x"90BF" when address_in = 16#21AF# else
		x"9508" when address_in = 16#21B0# else
		x"926F" when address_in = 16#21B1# else
		x"927F" when address_in = 16#21B2# else
		x"928F" when address_in = 16#21B3# else
		x"929F" when address_in = 16#21B4# else
		x"92AF" when address_in = 16#21B5# else
		x"92BF" when address_in = 16#21B6# else
		x"92DF" when address_in = 16#21B7# else
		x"92EF" when address_in = 16#21B8# else
		x"92FF" when address_in = 16#21B9# else
		x"930F" when address_in = 16#21BA# else
		x"931F" when address_in = 16#21BB# else
		x"93CF" when address_in = 16#21BC# else
		x"93DF" when address_in = 16#21BD# else
		x"2F08" when address_in = 16#21BE# else
		x"2F19" when address_in = 16#21BF# else
		x"2E86" when address_in = 16#21C0# else
		x"2E97" when address_in = 16#21C1# else
		x"2E64" when address_in = 16#21C2# else
		x"2E75" when address_in = 16#21C3# else
		x"B6DF" when address_in = 16#21C4# else
		x"94F8" when address_in = 16#21C5# else
		x"9180" when address_in = 16#21C6# else
		x"0102" when address_in = 16#21C7# else
		x"3084" when address_in = 16#21C8# else
		x"F411" when address_in = 16#21C9# else
		x"BEDF" when address_in = 16#21CA# else
		x"C05D" when address_in = 16#21CB# else
		x"E040" when address_in = 16#21CC# else
		x"24EE" when address_in = 16#21CD# else
		x"24FF" when address_in = 16#21CE# else
		x"2D3F" when address_in = 16#21CF# else
		x"2D2E" when address_in = 16#21D0# else
		x"2CAE" when address_in = 16#21D1# else
		x"2CBF" when address_in = 16#21D2# else
		x"2FF3" when address_in = 16#21D3# else
		x"2FE2" when address_in = 16#21D4# else
		x"0DEA" when address_in = 16#21D5# else
		x"1DFB" when address_in = 16#21D6# else
		x"5EE9" when address_in = 16#21D7# else
		x"4FFE" when address_in = 16#21D8# else
		x"8184" when address_in = 16#21D9# else
		x"8195" when address_in = 16#21DA# else
		x"2B89" when address_in = 16#21DB# else
		x"F009" when address_in = 16#21DC# else
		x"C03D" when address_in = 16#21DD# else
		x"E087" when address_in = 16#21DE# else
		x"E091" when address_in = 16#21DF# else
		x"940E" when address_in = 16#21E0# else
		x"241D" when address_in = 16#21E1# else
		x"3081" when address_in = 16#21E2# else
		x"F431" when address_in = 16#21E3# else
		x"E040" when address_in = 16#21E4# else
		x"2F60" when address_in = 16#21E5# else
		x"2F71" when address_in = 16#21E6# else
		x"2788" when address_in = 16#21E7# else
		x"2799" when address_in = 16#21E8# else
		x"C01A" when address_in = 16#21E9# else
		x"B781" when address_in = 16#21EA# else
		x"5F8F" when address_in = 16#21EB# else
		x"B722" when address_in = 16#21EC# else
		x"2799" when address_in = 16#21ED# else
		x"1B82" when address_in = 16#21EE# else
		x"0991" when address_in = 16#21EF# else
		x"1780" when address_in = 16#21F0# else
		x"0791" when address_in = 16#21F1# else
		x"F098" when address_in = 16#21F2# else
		x"E087" when address_in = 16#21F3# else
		x"E091" when address_in = 16#21F4# else
		x"940E" when address_in = 16#21F5# else
		x"241D" when address_in = 16#21F6# else
		x"2FA0" when address_in = 16#21F7# else
		x"2FB1" when address_in = 16#21F8# else
		x"27CC" when address_in = 16#21F9# else
		x"27DD" when address_in = 16#21FA# else
		x"3081" when address_in = 16#21FB# else
		x"F411" when address_in = 16#21FC# else
		x"E040" when address_in = 16#21FD# else
		x"C001" when address_in = 16#21FE# else
		x"E041" when address_in = 16#21FF# else
		x"2F6A" when address_in = 16#2200# else
		x"2F7B" when address_in = 16#2201# else
		x"2F8C" when address_in = 16#2202# else
		x"2F9D" when address_in = 16#2203# else
		x"940E" when address_in = 16#2204# else
		x"1D87" when address_in = 16#2205# else
		x"9180" when address_in = 16#2206# else
		x"0102" when address_in = 16#2207# else
		x"5F8F" when address_in = 16#2208# else
		x"9380" when address_in = 16#2209# else
		x"0102" when address_in = 16#220A# else
		x"2DFF" when address_in = 16#220B# else
		x"2DEE" when address_in = 16#220C# else
		x"0DEA" when address_in = 16#220D# else
		x"1DFB" when address_in = 16#220E# else
		x"5EE9" when address_in = 16#220F# else
		x"4FFE" when address_in = 16#2210# else
		x"8311" when address_in = 16#2211# else
		x"8300" when address_in = 16#2212# else
		x"8293" when address_in = 16#2213# else
		x"8282" when address_in = 16#2214# else
		x"8275" when address_in = 16#2215# else
		x"8264" when address_in = 16#2216# else
		x"BEDF" when address_in = 16#2217# else
		x"E080" when address_in = 16#2218# else
		x"E090" when address_in = 16#2219# else
		x"C010" when address_in = 16#221A# else
		x"5F4F" when address_in = 16#221B# else
		x"9408" when address_in = 16#221C# else
		x"1CA1" when address_in = 16#221D# else
		x"1CB1" when address_in = 16#221E# else
		x"5F2B" when address_in = 16#221F# else
		x"4F3F" when address_in = 16#2220# else
		x"E085" when address_in = 16#2221# else
		x"E090" when address_in = 16#2222# else
		x"0EE8" when address_in = 16#2223# else
		x"1EF9" when address_in = 16#2224# else
		x"3044" when address_in = 16#2225# else
		x"F408" when address_in = 16#2226# else
		x"CFAB" when address_in = 16#2227# else
		x"BEDF" when address_in = 16#2228# else
		x"EF84" when address_in = 16#2229# else
		x"EF9F" when address_in = 16#222A# else
		x"91DF" when address_in = 16#222B# else
		x"91CF" when address_in = 16#222C# else
		x"911F" when address_in = 16#222D# else
		x"910F" when address_in = 16#222E# else
		x"90FF" when address_in = 16#222F# else
		x"90EF" when address_in = 16#2230# else
		x"90DF" when address_in = 16#2231# else
		x"90BF" when address_in = 16#2232# else
		x"90AF" when address_in = 16#2233# else
		x"909F" when address_in = 16#2234# else
		x"908F" when address_in = 16#2235# else
		x"907F" when address_in = 16#2236# else
		x"906F" when address_in = 16#2237# else
		x"9508" when address_in = 16#2238# else
		x"2FB9" when address_in = 16#2239# else
		x"2FA8" when address_in = 16#223A# else
		x"B76F" when address_in = 16#223B# else
		x"94F8" when address_in = 16#223C# else
		x"E070" when address_in = 16#223D# else
		x"E020" when address_in = 16#223E# else
		x"E030" when address_in = 16#223F# else
		x"2F53" when address_in = 16#2240# else
		x"2F42" when address_in = 16#2241# else
		x"2FF3" when address_in = 16#2242# else
		x"2FE2" when address_in = 16#2243# else
		x"0FE4" when address_in = 16#2244# else
		x"1FF5" when address_in = 16#2245# else
		x"5EE9" when address_in = 16#2246# else
		x"4FFE" when address_in = 16#2247# else
		x"8184" when address_in = 16#2248# else
		x"8195" when address_in = 16#2249# else
		x"178A" when address_in = 16#224A# else
		x"079B" when address_in = 16#224B# else
		x"F459" when address_in = 16#224C# else
		x"8215" when address_in = 16#224D# else
		x"8214" when address_in = 16#224E# else
		x"9180" when address_in = 16#224F# else
		x"0102" when address_in = 16#2250# else
		x"5081" when address_in = 16#2251# else
		x"9380" when address_in = 16#2252# else
		x"0102" when address_in = 16#2253# else
		x"BF6F" when address_in = 16#2254# else
		x"E080" when address_in = 16#2255# else
		x"E090" when address_in = 16#2256# else
		x"9508" when address_in = 16#2257# else
		x"5F7F" when address_in = 16#2258# else
		x"5F4F" when address_in = 16#2259# else
		x"4F5F" when address_in = 16#225A# else
		x"5F2B" when address_in = 16#225B# else
		x"4F3F" when address_in = 16#225C# else
		x"3074" when address_in = 16#225D# else
		x"F318" when address_in = 16#225E# else
		x"BF6F" when address_in = 16#225F# else
		x"EE8A" when address_in = 16#2260# else
		x"EF9F" when address_in = 16#2261# else
		x"9508" when address_in = 16#2262# else
		x"921F" when address_in = 16#2263# else
		x"920F" when address_in = 16#2264# else
		x"B60F" when address_in = 16#2265# else
		x"920F" when address_in = 16#2266# else
		x"2411" when address_in = 16#2267# else
		x"932F" when address_in = 16#2268# else
		x"933F" when address_in = 16#2269# else
		x"934F" when address_in = 16#226A# else
		x"935F" when address_in = 16#226B# else
		x"936F" when address_in = 16#226C# else
		x"937F" when address_in = 16#226D# else
		x"938F" when address_in = 16#226E# else
		x"939F" when address_in = 16#226F# else
		x"93AF" when address_in = 16#2270# else
		x"93BF" when address_in = 16#2271# else
		x"93CF" when address_in = 16#2272# else
		x"93DF" when address_in = 16#2273# else
		x"93EF" when address_in = 16#2274# else
		x"93FF" when address_in = 16#2275# else
		x"B781" when address_in = 16#2276# else
		x"5F8F" when address_in = 16#2277# else
		x"2FC8" when address_in = 16#2278# else
		x"27DD" when address_in = 16#2279# else
		x"9180" when address_in = 16#227A# else
		x"0103" when address_in = 16#227B# else
		x"9190" when address_in = 16#227C# else
		x"0104" when address_in = 16#227D# else
		x"91A0" when address_in = 16#227E# else
		x"0105" when address_in = 16#227F# else
		x"91B0" when address_in = 16#2280# else
		x"0106" when address_in = 16#2281# else
		x"0F8C" when address_in = 16#2282# else
		x"1D91" when address_in = 16#2283# else
		x"1DA1" when address_in = 16#2284# else
		x"1DB1" when address_in = 16#2285# else
		x"9380" when address_in = 16#2286# else
		x"0103" when address_in = 16#2287# else
		x"9390" when address_in = 16#2288# else
		x"0104" when address_in = 16#2289# else
		x"93A0" when address_in = 16#228A# else
		x"0105" when address_in = 16#228B# else
		x"93B0" when address_in = 16#228C# else
		x"0106" when address_in = 16#228D# else
		x"E96C" when address_in = 16#228E# else
		x"E270" when address_in = 16#228F# else
		x"E080" when address_in = 16#2290# else
		x"940E" when address_in = 16#2291# else
		x"0B1A" when address_in = 16#2292# else
		x"9180" when address_in = 16#2293# else
		x"0102" when address_in = 16#2294# else
		x"2388" when address_in = 16#2295# else
		x"F059" when address_in = 16#2296# else
		x"2F8C" when address_in = 16#2297# else
		x"940E" when address_in = 16#2298# else
		x"1CEC" when address_in = 16#2299# else
		x"27AA" when address_in = 16#229A# else
		x"27BB" when address_in = 16#229B# else
		x"2F68" when address_in = 16#229C# else
		x"2F79" when address_in = 16#229D# else
		x"2F8A" when address_in = 16#229E# else
		x"2F9B" when address_in = 16#229F# else
		x"940E" when address_in = 16#22A0# else
		x"1CCD" when address_in = 16#22A1# else
		x"91FF" when address_in = 16#22A2# else
		x"91EF" when address_in = 16#22A3# else
		x"91DF" when address_in = 16#22A4# else
		x"91CF" when address_in = 16#22A5# else
		x"91BF" when address_in = 16#22A6# else
		x"91AF" when address_in = 16#22A7# else
		x"919F" when address_in = 16#22A8# else
		x"918F" when address_in = 16#22A9# else
		x"917F" when address_in = 16#22AA# else
		x"916F" when address_in = 16#22AB# else
		x"915F" when address_in = 16#22AC# else
		x"914F" when address_in = 16#22AD# else
		x"913F" when address_in = 16#22AE# else
		x"912F" when address_in = 16#22AF# else
		x"900F" when address_in = 16#22B0# else
		x"BE0F" when address_in = 16#22B1# else
		x"900F" when address_in = 16#22B2# else
		x"901F" when address_in = 16#22B3# else
		x"9518" when address_in = 16#22B4# else
		x"9210" when address_in = 16#22B5# else
		x"0130" when address_in = 16#22B6# else
		x"9210" when address_in = 16#22B7# else
		x"012F" when address_in = 16#22B8# else
		x"E080" when address_in = 16#22B9# else
		x"E090" when address_in = 16#22BA# else
		x"9508" when address_in = 16#22BB# else
		x"931F" when address_in = 16#22BC# else
		x"93CF" when address_in = 16#22BD# else
		x"93DF" when address_in = 16#22BE# else
		x"2F16" when address_in = 16#22BF# else
		x"2FD5" when address_in = 16#22C0# else
		x"2FC4" when address_in = 16#22C1# else
		x"940E" when address_in = 16#22C2# else
		x"0B28" when address_in = 16#22C3# else
		x"839A" when address_in = 16#22C4# else
		x"8389" when address_in = 16#22C5# else
		x"2B89" when address_in = 16#22C6# else
		x"F419" when address_in = 16#22C7# else
		x"EF8D" when address_in = 16#22C8# else
		x"EF9F" when address_in = 16#22C9# else
		x"C01C" when address_in = 16#22CA# else
		x"8318" when address_in = 16#22CB# else
		x"821C" when address_in = 16#22CC# else
		x"821B" when address_in = 16#22CD# else
		x"9180" when address_in = 16#22CE# else
		x"012F" when address_in = 16#22CF# else
		x"9190" when address_in = 16#22D0# else
		x"0130" when address_in = 16#22D1# else
		x"9700" when address_in = 16#22D2# else
		x"F429" when address_in = 16#22D3# else
		x"93D0" when address_in = 16#22D4# else
		x"0130" when address_in = 16#22D5# else
		x"93C0" when address_in = 16#22D6# else
		x"012F" when address_in = 16#22D7# else
		x"C00C" when address_in = 16#22D8# else
		x"2FF9" when address_in = 16#22D9# else
		x"2FE8" when address_in = 16#22DA# else
		x"8183" when address_in = 16#22DB# else
		x"8194" when address_in = 16#22DC# else
		x"2B89" when address_in = 16#22DD# else
		x"F021" when address_in = 16#22DE# else
		x"8003" when address_in = 16#22DF# else
		x"81F4" when address_in = 16#22E0# else
		x"2DE0" when address_in = 16#22E1# else
		x"CFF8" when address_in = 16#22E2# else
		x"83D4" when address_in = 16#22E3# else
		x"83C3" when address_in = 16#22E4# else
		x"E080" when address_in = 16#22E5# else
		x"E090" when address_in = 16#22E6# else
		x"91DF" when address_in = 16#22E7# else
		x"91CF" when address_in = 16#22E8# else
		x"911F" when address_in = 16#22E9# else
		x"9508" when address_in = 16#22EA# else
		x"91E0" when address_in = 16#22EB# else
		x"012F" when address_in = 16#22EC# else
		x"91F0" when address_in = 16#22ED# else
		x"0130" when address_in = 16#22EE# else
		x"2FAE" when address_in = 16#22EF# else
		x"2FBF" when address_in = 16#22F0# else
		x"9730" when address_in = 16#22F1# else
		x"F0D1" when address_in = 16#22F2# else
		x"17E8" when address_in = 16#22F3# else
		x"07F9" when address_in = 16#22F4# else
		x"F489" when address_in = 16#22F5# else
		x"8183" when address_in = 16#22F6# else
		x"8194" when address_in = 16#22F7# else
		x"17EA" when address_in = 16#22F8# else
		x"07FB" when address_in = 16#22F9# else
		x"F429" when address_in = 16#22FA# else
		x"9390" when address_in = 16#22FB# else
		x"0130" when address_in = 16#22FC# else
		x"9380" when address_in = 16#22FD# else
		x"012F" when address_in = 16#22FE# else
		x"C004" when address_in = 16#22FF# else
		x"2FFB" when address_in = 16#2300# else
		x"2FEA" when address_in = 16#2301# else
		x"8394" when address_in = 16#2302# else
		x"8383" when address_in = 16#2303# else
		x"E080" when address_in = 16#2304# else
		x"E090" when address_in = 16#2305# else
		x"9508" when address_in = 16#2306# else
		x"2FAE" when address_in = 16#2307# else
		x"2FBF" when address_in = 16#2308# else
		x"8003" when address_in = 16#2309# else
		x"81F4" when address_in = 16#230A# else
		x"2DE0" when address_in = 16#230B# else
		x"CFE4" when address_in = 16#230C# else
		x"EE8A" when address_in = 16#230D# else
		x"EF9F" when address_in = 16#230E# else
		x"9508" when address_in = 16#230F# else
		x"92DF" when address_in = 16#2310# else
		x"92EF" when address_in = 16#2311# else
		x"92FF" when address_in = 16#2312# else
		x"930F" when address_in = 16#2313# else
		x"931F" when address_in = 16#2314# else
		x"93CF" when address_in = 16#2315# else
		x"93DF" when address_in = 16#2316# else
		x"2EE8" when address_in = 16#2317# else
		x"2EF9" when address_in = 16#2318# else
		x"9140" when address_in = 16#2319# else
		x"012F" when address_in = 16#231A# else
		x"9150" when address_in = 16#231B# else
		x"0130" when address_in = 16#231C# else
		x"1541" when address_in = 16#231D# else
		x"0551" when address_in = 16#231E# else
		x"F409" when address_in = 16#231F# else
		x"C046" when address_in = 16#2320# else
		x"2FF9" when address_in = 16#2321# else
		x"2FE8" when address_in = 16#2322# else
		x"8124" when address_in = 16#2323# else
		x"8135" when address_in = 16#2324# else
		x"9180" when address_in = 16#2325# else
		x"0062" when address_in = 16#2326# else
		x"9190" when address_in = 16#2327# else
		x"0063" when address_in = 16#2328# else
		x"1728" when address_in = 16#2329# else
		x"0739" when address_in = 16#232A# else
		x"F419" when address_in = 16#232B# else
		x"E064" when address_in = 16#232C# else
		x"2ED6" when address_in = 16#232D# else
		x"C002" when address_in = 16#232E# else
		x"E031" when address_in = 16#232F# else
		x"2ED3" when address_in = 16#2330# else
		x"2F04" when address_in = 16#2331# else
		x"2F15" when address_in = 16#2332# else
		x"2B45" when address_in = 16#2333# else
		x"F409" when address_in = 16#2334# else
		x"C031" when address_in = 16#2335# else
		x"2FF1" when address_in = 16#2336# else
		x"2FE0" when address_in = 16#2337# else
		x"8180" when address_in = 16#2338# else
		x"218D" when address_in = 16#2339# else
		x"F129" when address_in = 16#233A# else
		x"81C1" when address_in = 16#233B# else
		x"81D2" when address_in = 16#233C# else
		x"819C" when address_in = 16#233D# else
		x"2DFF" when address_in = 16#233E# else
		x"2DEE" when address_in = 16#233F# else
		x"8180" when address_in = 16#2340# else
		x"1798" when address_in = 16#2341# else
		x"F0E9" when address_in = 16#2342# else
		x"818A" when address_in = 16#2343# else
		x"819B" when address_in = 16#2344# else
		x"27AA" when address_in = 16#2345# else
		x"27BB" when address_in = 16#2346# else
		x"0F88" when address_in = 16#2347# else
		x"1F99" when address_in = 16#2348# else
		x"1FAA" when address_in = 16#2349# else
		x"1FBB" when address_in = 16#234A# else
		x"960C" when address_in = 16#234B# else
		x"1DA1" when address_in = 16#234C# else
		x"1DB1" when address_in = 16#234D# else
		x"BFAB" when address_in = 16#234E# else
		x"2FF9" when address_in = 16#234F# else
		x"2FE8" when address_in = 16#2350# else
		x"95D8" when address_in = 16#2351# else
		x"2D20" when address_in = 16#2352# else
		x"B60B" when address_in = 16#2353# else
		x"9631" when address_in = 16#2354# else
		x"1C01" when address_in = 16#2355# else
		x"BE0B" when address_in = 16#2356# else
		x"95D8" when address_in = 16#2357# else
		x"2D30" when address_in = 16#2358# else
		x"2D7F" when address_in = 16#2359# else
		x"2D6E" when address_in = 16#235A# else
		x"818E" when address_in = 16#235B# else
		x"819F" when address_in = 16#235C# else
		x"2FE2" when address_in = 16#235D# else
		x"2FF3" when address_in = 16#235E# else
		x"9509" when address_in = 16#235F# else
		x"2FF1" when address_in = 16#2360# else
		x"2FE0" when address_in = 16#2361# else
		x"8103" when address_in = 16#2362# else
		x"8114" when address_in = 16#2363# else
		x"1501" when address_in = 16#2364# else
		x"0511" when address_in = 16#2365# else
		x"F679" when address_in = 16#2366# else
		x"91DF" when address_in = 16#2367# else
		x"91CF" when address_in = 16#2368# else
		x"911F" when address_in = 16#2369# else
		x"910F" when address_in = 16#236A# else
		x"90FF" when address_in = 16#236B# else
		x"90EF" when address_in = 16#236C# else
		x"90DF" when address_in = 16#236D# else
		x"9508" when address_in = 16#236E# else
		x"92EF" when address_in = 16#236F# else
		x"92FF" when address_in = 16#2370# else
		x"930F" when address_in = 16#2371# else
		x"931F" when address_in = 16#2372# else
		x"93CF" when address_in = 16#2373# else
		x"93DF" when address_in = 16#2374# else
		x"2EE8" when address_in = 16#2375# else
		x"2EF9" when address_in = 16#2376# else
		x"9180" when address_in = 16#2377# else
		x"012F" when address_in = 16#2378# else
		x"9190" when address_in = 16#2379# else
		x"0130" when address_in = 16#237A# else
		x"9700" when address_in = 16#237B# else
		x"F409" when address_in = 16#237C# else
		x"C033" when address_in = 16#237D# else
		x"2F08" when address_in = 16#237E# else
		x"2F19" when address_in = 16#237F# else
		x"2FF1" when address_in = 16#2380# else
		x"2FE0" when address_in = 16#2381# else
		x"8180" when address_in = 16#2382# else
		x"FF81" when address_in = 16#2383# else
		x"C025" when address_in = 16#2384# else
		x"81C1" when address_in = 16#2385# else
		x"81D2" when address_in = 16#2386# else
		x"819C" when address_in = 16#2387# else
		x"2DFF" when address_in = 16#2388# else
		x"2DEE" when address_in = 16#2389# else
		x"8181" when address_in = 16#238A# else
		x"1798" when address_in = 16#238B# else
		x"F0E9" when address_in = 16#238C# else
		x"818A" when address_in = 16#238D# else
		x"819B" when address_in = 16#238E# else
		x"27AA" when address_in = 16#238F# else
		x"27BB" when address_in = 16#2390# else
		x"0F88" when address_in = 16#2391# else
		x"1F99" when address_in = 16#2392# else
		x"1FAA" when address_in = 16#2393# else
		x"1FBB" when address_in = 16#2394# else
		x"960C" when address_in = 16#2395# else
		x"1DA1" when address_in = 16#2396# else
		x"1DB1" when address_in = 16#2397# else
		x"BFAB" when address_in = 16#2398# else
		x"2FF9" when address_in = 16#2399# else
		x"2FE8" when address_in = 16#239A# else
		x"95D8" when address_in = 16#239B# else
		x"2D20" when address_in = 16#239C# else
		x"B60B" when address_in = 16#239D# else
		x"9631" when address_in = 16#239E# else
		x"1C01" when address_in = 16#239F# else
		x"BE0B" when address_in = 16#23A0# else
		x"95D8" when address_in = 16#23A1# else
		x"2D30" when address_in = 16#23A2# else
		x"2D7F" when address_in = 16#23A3# else
		x"2D6E" when address_in = 16#23A4# else
		x"818E" when address_in = 16#23A5# else
		x"819F" when address_in = 16#23A6# else
		x"2FE2" when address_in = 16#23A7# else
		x"2FF3" when address_in = 16#23A8# else
		x"9509" when address_in = 16#23A9# else
		x"2FF1" when address_in = 16#23AA# else
		x"2FE0" when address_in = 16#23AB# else
		x"8103" when address_in = 16#23AC# else
		x"8114" when address_in = 16#23AD# else
		x"1501" when address_in = 16#23AE# else
		x"0511" when address_in = 16#23AF# else
		x"F679" when address_in = 16#23B0# else
		x"91DF" when address_in = 16#23B1# else
		x"91CF" when address_in = 16#23B2# else
		x"911F" when address_in = 16#23B3# else
		x"910F" when address_in = 16#23B4# else
		x"90FF" when address_in = 16#23B5# else
		x"90EF" when address_in = 16#23B6# else
		x"9508" when address_in = 16#23B7# else
		x"93CF" when address_in = 16#23B8# else
		x"93DF" when address_in = 16#23B9# else
		x"2FB7" when address_in = 16#23BA# else
		x"2FA6" when address_in = 16#23BB# else
		x"938D" when address_in = 16#23BC# else
		x"939C" when address_in = 16#23BD# else
		x"2FD9" when address_in = 16#23BE# else
		x"2FC8" when address_in = 16#23BF# else
		x"818A" when address_in = 16#23C0# else
		x"819B" when address_in = 16#23C1# else
		x"2FF7" when address_in = 16#23C2# else
		x"2FE6" when address_in = 16#23C3# else
		x"8393" when address_in = 16#23C4# else
		x"8382" when address_in = 16#23C5# else
		x"81EA" when address_in = 16#23C6# else
		x"81FB" when address_in = 16#23C7# else
		x"8371" when address_in = 16#23C8# else
		x"8360" when address_in = 16#23C9# else
		x"837B" when address_in = 16#23CA# else
		x"836A" when address_in = 16#23CB# else
		x"91DF" when address_in = 16#23CC# else
		x"91CF" when address_in = 16#23CD# else
		x"9508" when address_in = 16#23CE# else
		x"2FF9" when address_in = 16#23CF# else
		x"2FE8" when address_in = 16#23D0# else
		x"8180" when address_in = 16#23D1# else
		x"8191" when address_in = 16#23D2# else
		x"940E" when address_in = 16#23D3# else
		x"23B8" when address_in = 16#23D4# else
		x"9508" when address_in = 16#23D5# else
		x"940E" when address_in = 16#23D6# else
		x"23B8" when address_in = 16#23D7# else
		x"9508" when address_in = 16#23D8# else
		x"93CF" when address_in = 16#23D9# else
		x"93DF" when address_in = 16#23DA# else
		x"2FF9" when address_in = 16#23DB# else
		x"2FE8" when address_in = 16#23DC# else
		x"8142" when address_in = 16#23DD# else
		x"8153" when address_in = 16#23DE# else
		x"81A0" when address_in = 16#23DF# else
		x"81B1" when address_in = 16#23E0# else
		x"2FD5" when address_in = 16#23E1# else
		x"2FC4" when address_in = 16#23E2# else
		x"8128" when address_in = 16#23E3# else
		x"8139" when address_in = 16#23E4# else
		x"1728" when address_in = 16#23E5# else
		x"0739" when address_in = 16#23E6# else
		x"F039" when address_in = 16#23E7# else
		x"2FDB" when address_in = 16#23E8# else
		x"2FCA" when address_in = 16#23E9# else
		x"818A" when address_in = 16#23EA# else
		x"819B" when address_in = 16#23EB# else
		x"178E" when address_in = 16#23EC# else
		x"079F" when address_in = 16#23ED# else
		x"F491" when address_in = 16#23EE# else
		x"172E" when address_in = 16#23EF# else
		x"073F" when address_in = 16#23F0# else
		x"F499" when address_in = 16#23F1# else
		x"2FDB" when address_in = 16#23F2# else
		x"2FCA" when address_in = 16#23F3# else
		x"818A" when address_in = 16#23F4# else
		x"819B" when address_in = 16#23F5# else
		x"178E" when address_in = 16#23F6# else
		x"079F" when address_in = 16#23F7# else
		x"F461" when address_in = 16#23F8# else
		x"2FD5" when address_in = 16#23F9# else
		x"2FC4" when address_in = 16#23FA# else
		x"83B9" when address_in = 16#23FB# else
		x"83A8" when address_in = 16#23FC# else
		x"2FDB" when address_in = 16#23FD# else
		x"2FCA" when address_in = 16#23FE# else
		x"835B" when address_in = 16#23FF# else
		x"834A" when address_in = 16#2400# else
		x"8211" when address_in = 16#2401# else
		x"8210" when address_in = 16#2402# else
		x"8213" when address_in = 16#2403# else
		x"8212" when address_in = 16#2404# else
		x"91DF" when address_in = 16#2405# else
		x"91CF" when address_in = 16#2406# else
		x"9508" when address_in = 16#2407# else
		x"2FF9" when address_in = 16#2408# else
		x"2FE8" when address_in = 16#2409# else
		x"8180" when address_in = 16#240A# else
		x"8191" when address_in = 16#240B# else
		x"940E" when address_in = 16#240C# else
		x"23D9" when address_in = 16#240D# else
		x"9508" when address_in = 16#240E# else
		x"2FF9" when address_in = 16#240F# else
		x"2FE8" when address_in = 16#2410# else
		x"8182" when address_in = 16#2411# else
		x"8193" when address_in = 16#2412# else
		x"940E" when address_in = 16#2413# else
		x"23D9" when address_in = 16#2414# else
		x"9508" when address_in = 16#2415# else
		x"2FF9" when address_in = 16#2416# else
		x"2FE8" when address_in = 16#2417# else
		x"8393" when address_in = 16#2418# else
		x"8382" when address_in = 16#2419# else
		x"8391" when address_in = 16#241A# else
		x"8380" when address_in = 16#241B# else
		x"9508" when address_in = 16#241C# else
		x"2FF9" when address_in = 16#241D# else
		x"2FE8" when address_in = 16#241E# else
		x"E020" when address_in = 16#241F# else
		x"E030" when address_in = 16#2420# else
		x"8180" when address_in = 16#2421# else
		x"8191" when address_in = 16#2422# else
		x"178E" when address_in = 16#2423# else
		x"079F" when address_in = 16#2424# else
		x"F411" when address_in = 16#2425# else
		x"E021" when address_in = 16#2426# else
		x"E030" when address_in = 16#2427# else
		x"2F93" when address_in = 16#2428# else
		x"2F82" when address_in = 16#2429# else
		x"9508" when address_in = 16#242A# else
		x"E080" when address_in = 16#242B# else
		x"E090" when address_in = 16#242C# else
		x"9508" when address_in = 16#242D# else
		x"9390" when address_in = 16#242E# else
		x"0063" when address_in = 16#242F# else
		x"9380" when address_in = 16#2430# else
		x"0062" when address_in = 16#2431# else
		x"9508" when address_in = 16#2432# else
		x"9180" when address_in = 16#2433# else
		x"0062" when address_in = 16#2434# else
		x"9190" when address_in = 16#2435# else
		x"0063" when address_in = 16#2436# else
		x"9508" when address_in = 16#2437# else
		x"92AF" when address_in = 16#2438# else
		x"92BF" when address_in = 16#2439# else
		x"92CF" when address_in = 16#243A# else
		x"92DF" when address_in = 16#243B# else
		x"92EF" when address_in = 16#243C# else
		x"92FF" when address_in = 16#243D# else
		x"930F" when address_in = 16#243E# else
		x"931F" when address_in = 16#243F# else
		x"91E0" when address_in = 16#2440# else
		x"0077" when address_in = 16#2441# else
		x"9120" when address_in = 16#2442# else
		x"0070" when address_in = 16#2443# else
		x"9130" when address_in = 16#2444# else
		x"0071" when address_in = 16#2445# else
		x"9140" when address_in = 16#2446# else
		x"0072" when address_in = 16#2447# else
		x"9150" when address_in = 16#2448# else
		x"0073" when address_in = 16#2449# else
		x"9160" when address_in = 16#244A# else
		x"0074" when address_in = 16#244B# else
		x"9170" when address_in = 16#244C# else
		x"0075" when address_in = 16#244D# else
		x"9180" when address_in = 16#244E# else
		x"0076" when address_in = 16#244F# else
		x"2F9E" when address_in = 16#2450# else
		x"911F" when address_in = 16#2451# else
		x"910F" when address_in = 16#2452# else
		x"90FF" when address_in = 16#2453# else
		x"90EF" when address_in = 16#2454# else
		x"90DF" when address_in = 16#2455# else
		x"90CF" when address_in = 16#2456# else
		x"90BF" when address_in = 16#2457# else
		x"90AF" when address_in = 16#2458# else
		x"9508" when address_in = 16#2459# else
		x"93CF" when address_in = 16#245A# else
		x"93DF" when address_in = 16#245B# else
		x"2FF9" when address_in = 16#245C# else
		x"2FE8" when address_in = 16#245D# else
		x"E08C" when address_in = 16#245E# else
		x"E6A4" when address_in = 16#245F# else
		x"E0B0" when address_in = 16#2460# else
		x"2FCE" when address_in = 16#2461# else
		x"2FDF" when address_in = 16#2462# else
		x"900D" when address_in = 16#2463# else
		x"9209" when address_in = 16#2464# else
		x"958A" when address_in = 16#2465# else
		x"F7E1" when address_in = 16#2466# else
		x"2F8E" when address_in = 16#2467# else
		x"2F9F" when address_in = 16#2468# else
		x"91DF" when address_in = 16#2469# else
		x"91CF" when address_in = 16#246A# else
		x"9508" when address_in = 16#246B# else
		x"926F" when address_in = 16#246C# else
		x"927F" when address_in = 16#246D# else
		x"928F" when address_in = 16#246E# else
		x"929F" when address_in = 16#246F# else
		x"92AF" when address_in = 16#2470# else
		x"92BF" when address_in = 16#2471# else
		x"92CF" when address_in = 16#2472# else
		x"92DF" when address_in = 16#2473# else
		x"92EF" when address_in = 16#2474# else
		x"92FF" when address_in = 16#2475# else
		x"930F" when address_in = 16#2476# else
		x"931F" when address_in = 16#2477# else
		x"93CF" when address_in = 16#2478# else
		x"93DF" when address_in = 16#2479# else
		x"2E88" when address_in = 16#247A# else
		x"2E99" when address_in = 16#247B# else
		x"2FB9" when address_in = 16#247C# else
		x"2FA8" when address_in = 16#247D# else
		x"912D" when address_in = 16#247E# else
		x"913C" when address_in = 16#247F# else
		x"2FD7" when address_in = 16#2480# else
		x"2FC6" when address_in = 16#2481# else
		x"8188" when address_in = 16#2482# else
		x"8199" when address_in = 16#2483# else
		x"1728" when address_in = 16#2484# else
		x"0739" when address_in = 16#2485# else
		x"F029" when address_in = 16#2486# else
		x"EF2F" when address_in = 16#2487# else
		x"EF3F" when address_in = 16#2488# else
		x"EF4F" when address_in = 16#2489# else
		x"EF5F" when address_in = 16#248A# else
		x"C0B8" when address_in = 16#248B# else
		x"2DF9" when address_in = 16#248C# else
		x"2DE8" when address_in = 16#248D# else
		x"8182" when address_in = 16#248E# else
		x"8193" when address_in = 16#248F# else
		x"2FD7" when address_in = 16#2490# else
		x"2FC6" when address_in = 16#2491# else
		x"812A" when address_in = 16#2492# else
		x"813B" when address_in = 16#2493# else
		x"1B82" when address_in = 16#2494# else
		x"0B93" when address_in = 16#2495# else
		x"2FA8" when address_in = 16#2496# else
		x"2FB9" when address_in = 16#2497# else
		x"27CC" when address_in = 16#2498# else
		x"FDB7" when address_in = 16#2499# else
		x"95C0" when address_in = 16#249A# else
		x"2FDC" when address_in = 16#249B# else
		x"8184" when address_in = 16#249C# else
		x"8195" when address_in = 16#249D# else
		x"2FF7" when address_in = 16#249E# else
		x"2FE6" when address_in = 16#249F# else
		x"8124" when address_in = 16#24A0# else
		x"8135" when address_in = 16#24A1# else
		x"1B82" when address_in = 16#24A2# else
		x"0B93" when address_in = 16#24A3# else
		x"2EE8" when address_in = 16#24A4# else
		x"2EF9" when address_in = 16#24A5# else
		x"2700" when address_in = 16#24A6# else
		x"FCF7" when address_in = 16#24A7# else
		x"9500" when address_in = 16#24A8# else
		x"2F10" when address_in = 16#24A9# else
		x"2DF9" when address_in = 16#24AA# else
		x"2DE8" when address_in = 16#24AB# else
		x"8186" when address_in = 16#24AC# else
		x"8197" when address_in = 16#24AD# else
		x"2FF7" when address_in = 16#24AE# else
		x"2FE6" when address_in = 16#24AF# else
		x"8126" when address_in = 16#24B0# else
		x"8137" when address_in = 16#24B1# else
		x"1B82" when address_in = 16#24B2# else
		x"0B93" when address_in = 16#24B3# else
		x"2E68" when address_in = 16#24B4# else
		x"2E79" when address_in = 16#24B5# else
		x"2488" when address_in = 16#24B6# else
		x"FC77" when address_in = 16#24B7# else
		x"9480" when address_in = 16#24B8# else
		x"2C98" when address_in = 16#24B9# else
		x"30A0" when address_in = 16#24BA# else
		x"ECF0" when address_in = 16#24BB# else
		x"07BF" when address_in = 16#24BC# else
		x"EFFF" when address_in = 16#24BD# else
		x"07CF" when address_in = 16#24BE# else
		x"EFFF" when address_in = 16#24BF# else
		x"07DF" when address_in = 16#24C0# else
		x"F424" when address_in = 16#24C1# else
		x"E0A0" when address_in = 16#24C2# else
		x"ECB0" when address_in = 16#24C3# else
		x"EFCF" when address_in = 16#24C4# else
		x"EFDF" when address_in = 16#24C5# else
		x"E080" when address_in = 16#24C6# else
		x"16E8" when address_in = 16#24C7# else
		x"EC80" when address_in = 16#24C8# else
		x"06F8" when address_in = 16#24C9# else
		x"EF8F" when address_in = 16#24CA# else
		x"0708" when address_in = 16#24CB# else
		x"EF8F" when address_in = 16#24CC# else
		x"0718" when address_in = 16#24CD# else
		x"F43C" when address_in = 16#24CE# else
		x"2CE1" when address_in = 16#24CF# else
		x"EC30" when address_in = 16#24D0# else
		x"2EF3" when address_in = 16#24D1# else
		x"EF3F" when address_in = 16#24D2# else
		x"2F03" when address_in = 16#24D3# else
		x"EF3F" when address_in = 16#24D4# else
		x"2F13" when address_in = 16#24D5# else
		x"E0E0" when address_in = 16#24D6# else
		x"166E" when address_in = 16#24D7# else
		x"ECE0" when address_in = 16#24D8# else
		x"067E" when address_in = 16#24D9# else
		x"EFEF" when address_in = 16#24DA# else
		x"068E" when address_in = 16#24DB# else
		x"EFEF" when address_in = 16#24DC# else
		x"069E" when address_in = 16#24DD# else
		x"F43C" when address_in = 16#24DE# else
		x"2C61" when address_in = 16#24DF# else
		x"EC20" when address_in = 16#24E0# else
		x"2E72" when address_in = 16#24E1# else
		x"EF2F" when address_in = 16#24E2# else
		x"2E82" when address_in = 16#24E3# else
		x"EF2F" when address_in = 16#24E4# else
		x"2E92" when address_in = 16#24E5# else
		x"30A1" when address_in = 16#24E6# else
		x"E4F0" when address_in = 16#24E7# else
		x"07BF" when address_in = 16#24E8# else
		x"E0F0" when address_in = 16#24E9# else
		x"07CF" when address_in = 16#24EA# else
		x"E0F0" when address_in = 16#24EB# else
		x"07DF" when address_in = 16#24EC# else
		x"F024" when address_in = 16#24ED# else
		x"E0A0" when address_in = 16#24EE# else
		x"E4B0" when address_in = 16#24EF# else
		x"E0C0" when address_in = 16#24F0# else
		x"E0D0" when address_in = 16#24F1# else
		x"E081" when address_in = 16#24F2# else
		x"16E8" when address_in = 16#24F3# else
		x"E480" when address_in = 16#24F4# else
		x"06F8" when address_in = 16#24F5# else
		x"E080" when address_in = 16#24F6# else
		x"0708" when address_in = 16#24F7# else
		x"E080" when address_in = 16#24F8# else
		x"0718" when address_in = 16#24F9# else
		x"F02C" when address_in = 16#24FA# else
		x"2CE1" when address_in = 16#24FB# else
		x"E490" when address_in = 16#24FC# else
		x"2EF9" when address_in = 16#24FD# else
		x"2D01" when address_in = 16#24FE# else
		x"2D11" when address_in = 16#24FF# else
		x"E0E1" when address_in = 16#2500# else
		x"166E" when address_in = 16#2501# else
		x"E4E0" when address_in = 16#2502# else
		x"067E" when address_in = 16#2503# else
		x"E0E0" when address_in = 16#2504# else
		x"068E" when address_in = 16#2505# else
		x"E0E0" when address_in = 16#2506# else
		x"069E" when address_in = 16#2507# else
		x"F02C" when address_in = 16#2508# else
		x"2C61" when address_in = 16#2509# else
		x"E480" when address_in = 16#250A# else
		x"2E78" when address_in = 16#250B# else
		x"2C81" when address_in = 16#250C# else
		x"2C91" when address_in = 16#250D# else
		x"2F2A" when address_in = 16#250E# else
		x"2F3B" when address_in = 16#250F# else
		x"2F4C" when address_in = 16#2510# else
		x"2F5D" when address_in = 16#2511# else
		x"2F6A" when address_in = 16#2512# else
		x"2F7B" when address_in = 16#2513# else
		x"2F8C" when address_in = 16#2514# else
		x"2F9D" when address_in = 16#2515# else
		x"940E" when address_in = 16#2516# else
		x"2E88" when address_in = 16#2517# else
		x"2EA6" when address_in = 16#2518# else
		x"2EB7" when address_in = 16#2519# else
		x"2EC8" when address_in = 16#251A# else
		x"2ED9" when address_in = 16#251B# else
		x"2F51" when address_in = 16#251C# else
		x"2F40" when address_in = 16#251D# else
		x"2D3F" when address_in = 16#251E# else
		x"2D2E" when address_in = 16#251F# else
		x"2F91" when address_in = 16#2520# else
		x"2F80" when address_in = 16#2521# else
		x"2D7F" when address_in = 16#2522# else
		x"2D6E" when address_in = 16#2523# else
		x"940E" when address_in = 16#2524# else
		x"2E88" when address_in = 16#2525# else
		x"2EE6" when address_in = 16#2526# else
		x"2EF7" when address_in = 16#2527# else
		x"2F08" when address_in = 16#2528# else
		x"2F19" when address_in = 16#2529# else
		x"2D59" when address_in = 16#252A# else
		x"2D48" when address_in = 16#252B# else
		x"2D37" when address_in = 16#252C# else
		x"2D26" when address_in = 16#252D# else
		x"2D99" when address_in = 16#252E# else
		x"2D88" when address_in = 16#252F# else
		x"2D77" when address_in = 16#2530# else
		x"2D66" when address_in = 16#2531# else
		x"940E" when address_in = 16#2532# else
		x"2E88" when address_in = 16#2533# else
		x"2FB9" when address_in = 16#2534# else
		x"2FA8" when address_in = 16#2535# else
		x"2F97" when address_in = 16#2536# else
		x"2F86" when address_in = 16#2537# else
		x"2D5D" when address_in = 16#2538# else
		x"2D4C" when address_in = 16#2539# else
		x"2D3B" when address_in = 16#253A# else
		x"2D2A" when address_in = 16#253B# else
		x"0D2E" when address_in = 16#253C# else
		x"1D3F" when address_in = 16#253D# else
		x"1F40" when address_in = 16#253E# else
		x"1F51" when address_in = 16#253F# else
		x"0F28" when address_in = 16#2540# else
		x"1F39" when address_in = 16#2541# else
		x"1F4A" when address_in = 16#2542# else
		x"1F5B" when address_in = 16#2543# else
		x"2F95" when address_in = 16#2544# else
		x"2F84" when address_in = 16#2545# else
		x"2F73" when address_in = 16#2546# else
		x"2F62" when address_in = 16#2547# else
		x"91DF" when address_in = 16#2548# else
		x"91CF" when address_in = 16#2549# else
		x"911F" when address_in = 16#254A# else
		x"910F" when address_in = 16#254B# else
		x"90FF" when address_in = 16#254C# else
		x"90EF" when address_in = 16#254D# else
		x"90DF" when address_in = 16#254E# else
		x"90CF" when address_in = 16#254F# else
		x"90BF" when address_in = 16#2550# else
		x"90AF" when address_in = 16#2551# else
		x"909F" when address_in = 16#2552# else
		x"908F" when address_in = 16#2553# else
		x"907F" when address_in = 16#2554# else
		x"906F" when address_in = 16#2555# else
		x"9508" when address_in = 16#2556# else
		x"EF8D" when address_in = 16#2557# else
		x"EF9F" when address_in = 16#2558# else
		x"9508" when address_in = 16#2559# else
		x"E081" when address_in = 16#255A# else
		x"E090" when address_in = 16#255B# else
		x"9508" when address_in = 16#255C# else
		x"9180" when address_in = 16#255D# else
		x"0060" when address_in = 16#255E# else
		x"2799" when address_in = 16#255F# else
		x"9508" when address_in = 16#2560# else
		x"9180" when address_in = 16#2561# else
		x"0061" when address_in = 16#2562# else
		x"2799" when address_in = 16#2563# else
		x"9508" when address_in = 16#2564# else
		x"9380" when address_in = 16#2565# else
		x"0061" when address_in = 16#2566# else
		x"9508" when address_in = 16#2567# else
		x"B74F" when address_in = 16#2568# else
		x"94F8" when address_in = 16#2569# else
		x"9120" when address_in = 16#256A# else
		x"0062" when address_in = 16#256B# else
		x"9130" when address_in = 16#256C# else
		x"0063" when address_in = 16#256D# else
		x"2F93" when address_in = 16#256E# else
		x"2F82" when address_in = 16#256F# else
		x"E561" when address_in = 16#2570# else
		x"E377" when address_in = 16#2571# else
		x"940E" when address_in = 16#2572# else
		x"2E76" when address_in = 16#2573# else
		x"5A8F" when address_in = 16#2574# else
		x"4C98" when address_in = 16#2575# else
		x"9390" when address_in = 16#2576# else
		x"0132" when address_in = 16#2577# else
		x"9380" when address_in = 16#2578# else
		x"0131" when address_in = 16#2579# else
		x"9390" when address_in = 16#257A# else
		x"0134" when address_in = 16#257B# else
		x"9380" when address_in = 16#257C# else
		x"0133" when address_in = 16#257D# else
		x"2F93" when address_in = 16#257E# else
		x"2F82" when address_in = 16#257F# else
		x"E865" when address_in = 16#2580# else
		x"E07F" when address_in = 16#2581# else
		x"940E" when address_in = 16#2582# else
		x"2E76" when address_in = 16#2583# else
		x"578B" when address_in = 16#2584# else
		x"4F90" when address_in = 16#2585# else
		x"9390" when address_in = 16#2586# else
		x"0136" when address_in = 16#2587# else
		x"9380" when address_in = 16#2588# else
		x"0135" when address_in = 16#2589# else
		x"BF4F" when address_in = 16#258A# else
		x"9508" when address_in = 16#258B# else
		x"B78F" when address_in = 16#258C# else
		x"94F8" when address_in = 16#258D# else
		x"9120" when address_in = 16#258E# else
		x"0131" when address_in = 16#258F# else
		x"9130" when address_in = 16#2590# else
		x"0132" when address_in = 16#2591# else
		x"BF8F" when address_in = 16#2592# else
		x"2F83" when address_in = 16#2593# else
		x"1F88" when address_in = 16#2594# else
		x"2788" when address_in = 16#2595# else
		x"1F88" when address_in = 16#2596# else
		x"0F22" when address_in = 16#2597# else
		x"1F33" when address_in = 16#2598# else
		x"2388" when address_in = 16#2599# else
		x"F021" when address_in = 16#259A# else
		x"E08B" when address_in = 16#259B# else
		x"E190" when address_in = 16#259C# else
		x"2728" when address_in = 16#259D# else
		x"2739" when address_in = 16#259E# else
		x"5F2F" when address_in = 16#259F# else
		x"4F3F" when address_in = 16#25A0# else
		x"B78F" when address_in = 16#25A1# else
		x"94F8" when address_in = 16#25A2# else
		x"9330" when address_in = 16#25A3# else
		x"0132" when address_in = 16#25A4# else
		x"9320" when address_in = 16#25A5# else
		x"0131" when address_in = 16#25A6# else
		x"BF8F" when address_in = 16#25A7# else
		x"9180" when address_in = 16#25A8# else
		x"0135" when address_in = 16#25A9# else
		x"9190" when address_in = 16#25AA# else
		x"0136" when address_in = 16#25AB# else
		x"2782" when address_in = 16#25AC# else
		x"2793" when address_in = 16#25AD# else
		x"9508" when address_in = 16#25AE# else
		x"9210" when address_in = 16#25AF# else
		x"0147" when address_in = 16#25B0# else
		x"9210" when address_in = 16#25B1# else
		x"0149" when address_in = 16#25B2# else
		x"9210" when address_in = 16#25B3# else
		x"0148" when address_in = 16#25B4# else
		x"940E" when address_in = 16#25B5# else
		x"2433" when address_in = 16#25B6# else
		x"940E" when address_in = 16#25B7# else
		x"26CA" when address_in = 16#25B8# else
		x"E18C" when address_in = 16#25B9# else
		x"E099" when address_in = 16#25BA# else
		x"27AA" when address_in = 16#25BB# else
		x"FD97" when address_in = 16#25BC# else
		x"95A0" when address_in = 16#25BD# else
		x"2FBA" when address_in = 16#25BE# else
		x"95B6" when address_in = 16#25BF# else
		x"95A7" when address_in = 16#25C0# else
		x"9597" when address_in = 16#25C1# else
		x"9587" when address_in = 16#25C2# else
		x"940E" when address_in = 16#25C3# else
		x"0D10" when address_in = 16#25C4# else
		x"E387" when address_in = 16#25C5# else
		x"E091" when address_in = 16#25C6# else
		x"940E" when address_in = 16#25C7# else
		x"116D" when address_in = 16#25C8# else
		x"9508" when address_in = 16#25C9# else
		x"93CF" when address_in = 16#25CA# else
		x"93DF" when address_in = 16#25CB# else
		x"2FD9" when address_in = 16#25CC# else
		x"2FC8" when address_in = 16#25CD# else
		x"EC60" when address_in = 16#25CE# else
		x"E488" when address_in = 16#25CF# else
		x"940E" when address_in = 16#25D0# else
		x"2C68" when address_in = 16#25D1# else
		x"2388" when address_in = 16#25D2# else
		x"F021" when address_in = 16#25D3# else
		x"E488" when address_in = 16#25D4# else
		x"940E" when address_in = 16#25D5# else
		x"2C8E" when address_in = 16#25D6# else
		x"C00C" when address_in = 16#25D7# else
		x"E448" when address_in = 16#25D8# else
		x"816F" when address_in = 16#25D9# else
		x"2F8C" when address_in = 16#25DA# else
		x"2F9D" when address_in = 16#25DB# else
		x"940E" when address_in = 16#25DC# else
		x"2CD1" when address_in = 16#25DD# else
		x"2388" when address_in = 16#25DE# else
		x"F421" when address_in = 16#25DF# else
		x"E082" when address_in = 16#25E0# else
		x"9380" when address_in = 16#25E1# else
		x"0147" when address_in = 16#25E2# else
		x"C011" when address_in = 16#25E3# else
		x"E081" when address_in = 16#25E4# else
		x"9380" when address_in = 16#25E5# else
		x"0147" when address_in = 16#25E6# else
		x"2F6C" when address_in = 16#25E7# else
		x"2F7D" when address_in = 16#25E8# else
		x"E387" when address_in = 16#25E9# else
		x"E091" when address_in = 16#25EA# else
		x"940E" when address_in = 16#25EB# else
		x"1180" when address_in = 16#25EC# else
		x"E020" when address_in = 16#25ED# else
		x"E031" when address_in = 16#25EE# else
		x"E040" when address_in = 16#25EF# else
		x"E050" when address_in = 16#25F0# else
		x"E060" when address_in = 16#25F1# else
		x"E488" when address_in = 16#25F2# else
		x"940E" when address_in = 16#25F3# else
		x"1FCD" when address_in = 16#25F4# else
		x"91DF" when address_in = 16#25F5# else
		x"91CF" when address_in = 16#25F6# else
		x"9508" when address_in = 16#25F7# else
		x"931F" when address_in = 16#25F8# else
		x"93CF" when address_in = 16#25F9# else
		x"93DF" when address_in = 16#25FA# else
		x"2FD9" when address_in = 16#25FB# else
		x"2FC8" when address_in = 16#25FC# else
		x"858A" when address_in = 16#25FD# else
		x"859B" when address_in = 16#25FE# else
		x"FF82" when address_in = 16#25FF# else
		x"C00E" when address_in = 16#2600# else
		x"B184" when address_in = 16#2601# else
		x"2799" when address_in = 16#2602# else
		x"718E" when address_in = 16#2603# else
		x"7090" when address_in = 16#2604# else
		x"9595" when address_in = 16#2605# else
		x"9587" when address_in = 16#2606# else
		x"9595" when address_in = 16#2607# else
		x"9587" when address_in = 16#2608# else
		x"2F48" when address_in = 16#2609# else
		x"E468" when address_in = 16#260A# else
		x"8588" when address_in = 16#260B# else
		x"8599" when address_in = 16#260C# else
		x"940E" when address_in = 16#260D# else
		x"0700" when address_in = 16#260E# else
		x"B71F" when address_in = 16#260F# else
		x"94F8" when address_in = 16#2610# else
		x"9180" when address_in = 16#2611# else
		x"0147" when address_in = 16#2612# else
		x"2388" when address_in = 16#2613# else
		x"F449" when address_in = 16#2614# else
		x"93D0" when address_in = 16#2615# else
		x"0149" when address_in = 16#2616# else
		x"93C0" when address_in = 16#2617# else
		x"0148" when address_in = 16#2618# else
		x"2F8C" when address_in = 16#2619# else
		x"2F9D" when address_in = 16#261A# else
		x"940E" when address_in = 16#261B# else
		x"25CA" when address_in = 16#261C# else
		x"C006" when address_in = 16#261D# else
		x"2F6C" when address_in = 16#261E# else
		x"2F7D" when address_in = 16#261F# else
		x"E387" when address_in = 16#2620# else
		x"E091" when address_in = 16#2621# else
		x"940E" when address_in = 16#2622# else
		x"1180" when address_in = 16#2623# else
		x"BF1F" when address_in = 16#2624# else
		x"91DF" when address_in = 16#2625# else
		x"91CF" when address_in = 16#2626# else
		x"911F" when address_in = 16#2627# else
		x"9508" when address_in = 16#2628# else
		x"931F" when address_in = 16#2629# else
		x"93CF" when address_in = 16#262A# else
		x"93DF" when address_in = 16#262B# else
		x"2FF7" when address_in = 16#262C# else
		x"2FE6" when address_in = 16#262D# else
		x"B71F" when address_in = 16#262E# else
		x"94F8" when address_in = 16#262F# else
		x"8186" when address_in = 16#2630# else
		x"2799" when address_in = 16#2631# else
		x"3086" when address_in = 16#2632# else
		x"0591" when address_in = 16#2633# else
		x"F0C9" when address_in = 16#2634# else
		x"3087" when address_in = 16#2635# else
		x"0591" when address_in = 16#2636# else
		x"F434" when address_in = 16#2637# else
		x"9700" when address_in = 16#2638# else
		x"F061" when address_in = 16#2639# else
		x"9702" when address_in = 16#263A# else
		x"F409" when address_in = 16#263B# else
		x"C047" when address_in = 16#263C# else
		x"C074" when address_in = 16#263D# else
		x"308F" when address_in = 16#263E# else
		x"0591" when address_in = 16#263F# else
		x"F409" when address_in = 16#2640# else
		x"C055" when address_in = 16#2641# else
		x"3482" when address_in = 16#2642# else
		x"0591" when address_in = 16#2643# else
		x"F071" when address_in = 16#2644# else
		x"C06C" when address_in = 16#2645# else
		x"9210" when address_in = 16#2646# else
		x"0147" when address_in = 16#2647# else
		x"E041" when address_in = 16#2648# else
		x"E060" when address_in = 16#2649# else
		x"E488" when address_in = 16#264A# else
		x"940E" when address_in = 16#264B# else
		x"1F15" when address_in = 16#264C# else
		x"C068" when address_in = 16#264D# else
		x"E060" when address_in = 16#264E# else
		x"E488" when address_in = 16#264F# else
		x"940E" when address_in = 16#2650# else
		x"1EEF" when address_in = 16#2651# else
		x"C063" when address_in = 16#2652# else
		x"8582" when address_in = 16#2653# else
		x"9120" when address_in = 16#2654# else
		x"0148" when address_in = 16#2655# else
		x"9130" when address_in = 16#2656# else
		x"0149" when address_in = 16#2657# else
		x"9210" when address_in = 16#2658# else
		x"0149" when address_in = 16#2659# else
		x"9210" when address_in = 16#265A# else
		x"0148" when address_in = 16#265B# else
		x"E060" when address_in = 16#265C# else
		x"FF81" when address_in = 16#265D# else
		x"E061" when address_in = 16#265E# else
		x"E448" when address_in = 16#265F# else
		x"2F93" when address_in = 16#2660# else
		x"2F82" when address_in = 16#2661# else
		x"940E" when address_in = 16#2662# else
		x"13C4" when address_in = 16#2663# else
		x"E387" when address_in = 16#2664# else
		x"E091" when address_in = 16#2665# else
		x"940E" when address_in = 16#2666# else
		x"11CE" when address_in = 16#2667# else
		x"2FD9" when address_in = 16#2668# else
		x"2FC8" when address_in = 16#2669# else
		x"9390" when address_in = 16#266A# else
		x"0149" when address_in = 16#266B# else
		x"9380" when address_in = 16#266C# else
		x"0148" when address_in = 16#266D# else
		x"9700" when address_in = 16#266E# else
		x"F109" when address_in = 16#266F# else
		x"E448" when address_in = 16#2670# else
		x"816F" when address_in = 16#2671# else
		x"940E" when address_in = 16#2672# else
		x"2CD1" when address_in = 16#2673# else
		x"2388" when address_in = 16#2674# else
		x"F051" when address_in = 16#2675# else
		x"E081" when address_in = 16#2676# else
		x"9380" when address_in = 16#2677# else
		x"0147" when address_in = 16#2678# else
		x"2F6C" when address_in = 16#2679# else
		x"2F7D" when address_in = 16#267A# else
		x"E387" when address_in = 16#267B# else
		x"E091" when address_in = 16#267C# else
		x"940E" when address_in = 16#267D# else
		x"1180" when address_in = 16#267E# else
		x"C029" when address_in = 16#267F# else
		x"E082" when address_in = 16#2680# else
		x"9380" when address_in = 16#2681# else
		x"0147" when address_in = 16#2682# else
		x"C032" when address_in = 16#2683# else
		x"E387" when address_in = 16#2684# else
		x"E091" when address_in = 16#2685# else
		x"940E" when address_in = 16#2686# else
		x"11CE" when address_in = 16#2687# else
		x"9390" when address_in = 16#2688# else
		x"0149" when address_in = 16#2689# else
		x"9380" when address_in = 16#268A# else
		x"0148" when address_in = 16#268B# else
		x"9700" when address_in = 16#268C# else
		x"F019" when address_in = 16#268D# else
		x"940E" when address_in = 16#268E# else
		x"25CA" when address_in = 16#268F# else
		x"C025" when address_in = 16#2690# else
		x"E488" when address_in = 16#2691# else
		x"940E" when address_in = 16#2692# else
		x"2C8E" when address_in = 16#2693# else
		x"9210" when address_in = 16#2694# else
		x"0147" when address_in = 16#2695# else
		x"C01F" when address_in = 16#2696# else
		x"E488" when address_in = 16#2697# else
		x"940E" when address_in = 16#2698# else
		x"2C8E" when address_in = 16#2699# else
		x"9180" when address_in = 16#269A# else
		x"0148" when address_in = 16#269B# else
		x"9190" when address_in = 16#269C# else
		x"0149" when address_in = 16#269D# else
		x"9210" when address_in = 16#269E# else
		x"0149" when address_in = 16#269F# else
		x"9210" when address_in = 16#26A0# else
		x"0148" when address_in = 16#26A1# else
		x"E448" when address_in = 16#26A2# else
		x"E060" when address_in = 16#26A3# else
		x"940E" when address_in = 16#26A4# else
		x"13C4" when address_in = 16#26A5# else
		x"E081" when address_in = 16#26A6# else
		x"9380" when address_in = 16#26A7# else
		x"0147" when address_in = 16#26A8# else
		x"E020" when address_in = 16#26A9# else
		x"E031" when address_in = 16#26AA# else
		x"E040" when address_in = 16#26AB# else
		x"E050" when address_in = 16#26AC# else
		x"E060" when address_in = 16#26AD# else
		x"E488" when address_in = 16#26AE# else
		x"940E" when address_in = 16#26AF# else
		x"1FCD" when address_in = 16#26B0# else
		x"C004" when address_in = 16#26B1# else
		x"BF1F" when address_in = 16#26B2# else
		x"EE8A" when address_in = 16#26B3# else
		x"EF9F" when address_in = 16#26B4# else
		x"C003" when address_in = 16#26B5# else
		x"BF1F" when address_in = 16#26B6# else
		x"E080" when address_in = 16#26B7# else
		x"E090" when address_in = 16#26B8# else
		x"91DF" when address_in = 16#26B9# else
		x"91CF" when address_in = 16#26BA# else
		x"911F" when address_in = 16#26BB# else
		x"9508" when address_in = 16#26BC# else
		x"9120" when address_in = 16#26BD# else
		x"0078" when address_in = 16#26BE# else
		x"9130" when address_in = 16#26BF# else
		x"0079" when address_in = 16#26C0# else
		x"1782" when address_in = 16#26C1# else
		x"0793" when address_in = 16#26C2# else
		x"F019" when address_in = 16#26C3# else
		x"EE8A" when address_in = 16#26C4# else
		x"EF9F" when address_in = 16#26C5# else
		x"9508" when address_in = 16#26C6# else
		x"E080" when address_in = 16#26C7# else
		x"E090" when address_in = 16#26C8# else
		x"9508" when address_in = 16#26C9# else
		x"9390" when address_in = 16#26CA# else
		x"0079" when address_in = 16#26CB# else
		x"9380" when address_in = 16#26CC# else
		x"0078" when address_in = 16#26CD# else
		x"9508" when address_in = 16#26CE# else
		x"2799" when address_in = 16#26CF# else
		x"3085" when address_in = 16#26D0# else
		x"0591" when address_in = 16#26D1# else
		x"F131" when address_in = 16#26D2# else
		x"3086" when address_in = 16#26D3# else
		x"0591" when address_in = 16#26D4# else
		x"F47C" when address_in = 16#26D5# else
		x"3082" when address_in = 16#26D6# else
		x"0591" when address_in = 16#26D7# else
		x"F0D1" when address_in = 16#26D8# else
		x"3083" when address_in = 16#26D9# else
		x"0591" when address_in = 16#26DA# else
		x"F41C" when address_in = 16#26DB# else
		x"9701" when address_in = 16#26DC# else
		x"F099" when address_in = 16#26DD# else
		x"C028" when address_in = 16#26DE# else
		x"3083" when address_in = 16#26DF# else
		x"0591" when address_in = 16#26E0# else
		x"F099" when address_in = 16#26E1# else
		x"9704" when address_in = 16#26E2# else
		x"F099" when address_in = 16#26E3# else
		x"C022" when address_in = 16#26E4# else
		x"3087" when address_in = 16#26E5# else
		x"0591" when address_in = 16#26E6# else
		x"F0A9" when address_in = 16#26E7# else
		x"3087" when address_in = 16#26E8# else
		x"0591" when address_in = 16#26E9# else
		x"F084" when address_in = 16#26EA# else
		x"3088" when address_in = 16#26EB# else
		x"0591" when address_in = 16#26EC# else
		x"F091" when address_in = 16#26ED# else
		x"9709" when address_in = 16#26EE# else
		x"F099" when address_in = 16#26EF# else
		x"C016" when address_in = 16#26F0# else
		x"98DA" when address_in = 16#26F1# else
		x"C014" when address_in = 16#26F2# else
		x"98D9" when address_in = 16#26F3# else
		x"C012" when address_in = 16#26F4# else
		x"98D8" when address_in = 16#26F5# else
		x"C010" when address_in = 16#26F6# else
		x"9ADA" when address_in = 16#26F7# else
		x"C00E" when address_in = 16#26F8# else
		x"9AD9" when address_in = 16#26F9# else
		x"C00C" when address_in = 16#26FA# else
		x"9AD8" when address_in = 16#26FB# else
		x"C00A" when address_in = 16#26FC# else
		x"B38B" when address_in = 16#26FD# else
		x"E094" when address_in = 16#26FE# else
		x"C005" when address_in = 16#26FF# else
		x"B38B" when address_in = 16#2700# else
		x"E092" when address_in = 16#2701# else
		x"C002" when address_in = 16#2702# else
		x"B38B" when address_in = 16#2703# else
		x"E091" when address_in = 16#2704# else
		x"2789" when address_in = 16#2705# else
		x"BB8B" when address_in = 16#2706# else
		x"E080" when address_in = 16#2707# else
		x"E090" when address_in = 16#2708# else
		x"9508" when address_in = 16#2709# else
		x"9180" when address_in = 16#270A# else
		x"014A" when address_in = 16#270B# else
		x"2388" when address_in = 16#270C# else
		x"F451" when address_in = 16#270D# else
		x"B79F" when address_in = 16#270E# else
		x"94F8" when address_in = 16#270F# else
		x"E383" when address_in = 16#2710# else
		x"B989" when address_in = 16#2711# else
		x"E988" when address_in = 16#2712# else
		x"B98A" when address_in = 16#2713# else
		x"BF9F" when address_in = 16#2714# else
		x"E081" when address_in = 16#2715# else
		x"9380" when address_in = 16#2716# else
		x"014A" when address_in = 16#2717# else
		x"E080" when address_in = 16#2718# else
		x"E090" when address_in = 16#2719# else
		x"9508" when address_in = 16#271A# else
		x"E080" when address_in = 16#271B# else
		x"9380" when address_in = 16#271C# else
		x"014F" when address_in = 16#271D# else
		x"9380" when address_in = 16#271E# else
		x"015B" when address_in = 16#271F# else
		x"940E" when address_in = 16#2720# else
		x"270A" when address_in = 16#2721# else
		x"E091" when address_in = 16#2722# else
		x"E4EF" when address_in = 16#2723# else
		x"E0F1" when address_in = 16#2724# else
		x"2F89" when address_in = 16#2725# else
		x"8214" when address_in = 16#2726# else
		x"8213" when address_in = 16#2727# else
		x"8610" when address_in = 16#2728# else
		x"8217" when address_in = 16#2729# else
		x"8216" when address_in = 16#272A# else
		x"8215" when address_in = 16#272B# else
		x"8612" when address_in = 16#272C# else
		x"8613" when address_in = 16#272D# else
		x"8211" when address_in = 16#272E# else
		x"8212" when address_in = 16#272F# else
		x"8390" when address_in = 16#2730# else
		x"5081" when address_in = 16#2731# else
		x"963C" when address_in = 16#2732# else
		x"FF87" when address_in = 16#2733# else
		x"CFF1" when address_in = 16#2734# else
		x"9508" when address_in = 16#2735# else
		x"FF86" when address_in = 16#2736# else
		x"C004" when address_in = 16#2737# else
		x"9180" when address_in = 16#2738# else
		x"014F" when address_in = 16#2739# else
		x"2799" when address_in = 16#273A# else
		x"9508" when address_in = 16#273B# else
		x"9180" when address_in = 16#273C# else
		x"015B" when address_in = 16#273D# else
		x"2799" when address_in = 16#273E# else
		x"9508" when address_in = 16#273F# else
		x"2FF9" when address_in = 16#2740# else
		x"2FE8" when address_in = 16#2741# else
		x"9180" when address_in = 16#2742# else
		x"014F" when address_in = 16#2743# else
		x"3081" when address_in = 16#2744# else
		x"F019" when address_in = 16#2745# else
		x"EF80" when address_in = 16#2746# else
		x"EF9F" when address_in = 16#2747# else
		x"9508" when address_in = 16#2748# else
		x"2F84" when address_in = 16#2749# else
		x"7D81" when address_in = 16#274A# else
		x"9380" when address_in = 16#274B# else
		x"015A" when address_in = 16#274C# else
		x"FF87" when address_in = 16#274D# else
		x"C00E" when address_in = 16#274E# else
		x"93F0" when address_in = 16#274F# else
		x"0153" when address_in = 16#2750# else
		x"93E0" when address_in = 16#2751# else
		x"0152" when address_in = 16#2752# else
		x"8187" when address_in = 16#2753# else
		x"9380" when address_in = 16#2754# else
		x"0158" when address_in = 16#2755# else
		x"8580" when address_in = 16#2756# else
		x"8591" when address_in = 16#2757# else
		x"9390" when address_in = 16#2758# else
		x"0155" when address_in = 16#2759# else
		x"9380" when address_in = 16#275A# else
		x"0154" when address_in = 16#275B# else
		x"C006" when address_in = 16#275C# else
		x"93F0" when address_in = 16#275D# else
		x"0155" when address_in = 16#275E# else
		x"93E0" when address_in = 16#275F# else
		x"0154" when address_in = 16#2760# else
		x"9360" when address_in = 16#2761# else
		x"0158" when address_in = 16#2762# else
		x"9210" when address_in = 16#2763# else
		x"0159" when address_in = 16#2764# else
		x"E082" when address_in = 16#2765# else
		x"9380" when address_in = 16#2766# else
		x"014F" when address_in = 16#2767# else
		x"E081" when address_in = 16#2768# else
		x"9380" when address_in = 16#2769# else
		x"0151" when address_in = 16#276A# else
		x"9A56" when address_in = 16#276B# else
		x"E78E" when address_in = 16#276C# else
		x"B98C" when address_in = 16#276D# else
		x"E080" when address_in = 16#276E# else
		x"E090" when address_in = 16#276F# else
		x"9508" when address_in = 16#2770# else
		x"93CF" when address_in = 16#2771# else
		x"2FC8" when address_in = 16#2772# else
		x"9180" when address_in = 16#2773# else
		x"015B" when address_in = 16#2774# else
		x"3081" when address_in = 16#2775# else
		x"F019" when address_in = 16#2776# else
		x"EF80" when address_in = 16#2777# else
		x"EF9F" when address_in = 16#2778# else
		x"C035" when address_in = 16#2779# else
		x"2F86" when address_in = 16#277A# else
		x"7D81" when address_in = 16#277B# else
		x"9380" when address_in = 16#277C# else
		x"0166" when address_in = 16#277D# else
		x"FF67" when address_in = 16#277E# else
		x"C007" when address_in = 16#277F# else
		x"940E" when address_in = 16#2780# else
		x"12DE" when address_in = 16#2781# else
		x"9390" when address_in = 16#2782# else
		x"015F" when address_in = 16#2783# else
		x"9380" when address_in = 16#2784# else
		x"015E" when address_in = 16#2785# else
		x"C012" when address_in = 16#2786# else
		x"B184" when address_in = 16#2787# else
		x"2799" when address_in = 16#2788# else
		x"718E" when address_in = 16#2789# else
		x"7090" when address_in = 16#278A# else
		x"9595" when address_in = 16#278B# else
		x"9587" when address_in = 16#278C# else
		x"9595" when address_in = 16#278D# else
		x"9587" when address_in = 16#278E# else
		x"2F48" when address_in = 16#278F# else
		x"E462" when address_in = 16#2790# else
		x"2F8C" when address_in = 16#2791# else
		x"2799" when address_in = 16#2792# else
		x"940E" when address_in = 16#2793# else
		x"0889" when address_in = 16#2794# else
		x"9390" when address_in = 16#2795# else
		x"0161" when address_in = 16#2796# else
		x"9380" when address_in = 16#2797# else
		x"0160" when address_in = 16#2798# else
		x"2B89" when address_in = 16#2799# else
		x"F419" when address_in = 16#279A# else
		x"EF84" when address_in = 16#279B# else
		x"EF9F" when address_in = 16#279C# else
		x"C011" when address_in = 16#279D# else
		x"93C0" when address_in = 16#279E# else
		x"0164" when address_in = 16#279F# else
		x"9210" when address_in = 16#27A0# else
		x"0165" when address_in = 16#27A1# else
		x"9210" when address_in = 16#27A2# else
		x"0163" when address_in = 16#27A3# else
		x"9210" when address_in = 16#27A4# else
		x"0162" when address_in = 16#27A5# else
		x"E082" when address_in = 16#27A6# else
		x"9380" when address_in = 16#27A7# else
		x"015B" when address_in = 16#27A8# else
		x"E081" when address_in = 16#27A9# else
		x"9380" when address_in = 16#27AA# else
		x"015D" when address_in = 16#27AB# else
		x"9A57" when address_in = 16#27AC# else
		x"E080" when address_in = 16#27AD# else
		x"E090" when address_in = 16#27AE# else
		x"91CF" when address_in = 16#27AF# else
		x"9508" when address_in = 16#27B0# else
		x"9140" when address_in = 16#27B1# else
		x"0166" when address_in = 16#27B2# else
		x"2F84" when address_in = 16#27B3# else
		x"2799" when address_in = 16#27B4# else
		x"2F28" when address_in = 16#27B5# else
		x"2F39" when address_in = 16#27B6# else
		x"7220" when address_in = 16#27B7# else
		x"7030" when address_in = 16#27B8# else
		x"FF85" when address_in = 16#27B9# else
		x"C014" when address_in = 16#27BA# else
		x"B78F" when address_in = 16#27BB# else
		x"94F8" when address_in = 16#27BC# else
		x"7D4F" when address_in = 16#27BD# else
		x"9340" when address_in = 16#27BE# else
		x"0166" when address_in = 16#27BF# else
		x"BF8F" when address_in = 16#27C0# else
		x"9180" when address_in = 16#27C1# else
		x"0166" when address_in = 16#27C2# else
		x"FF87" when address_in = 16#27C3# else
		x"C005" when address_in = 16#27C4# else
		x"9180" when address_in = 16#27C5# else
		x"015E" when address_in = 16#27C6# else
		x"9190" when address_in = 16#27C7# else
		x"015F" when address_in = 16#27C8# else
		x"9508" when address_in = 16#27C9# else
		x"9180" when address_in = 16#27CA# else
		x"0160" when address_in = 16#27CB# else
		x"9190" when address_in = 16#27CC# else
		x"0161" when address_in = 16#27CD# else
		x"9508" when address_in = 16#27CE# else
		x"2F93" when address_in = 16#27CF# else
		x"2F82" when address_in = 16#27D0# else
		x"9508" when address_in = 16#27D1# else
		x"921F" when address_in = 16#27D2# else
		x"920F" when address_in = 16#27D3# else
		x"B60F" when address_in = 16#27D4# else
		x"920F" when address_in = 16#27D5# else
		x"2411" when address_in = 16#27D6# else
		x"932F" when address_in = 16#27D7# else
		x"933F" when address_in = 16#27D8# else
		x"934F" when address_in = 16#27D9# else
		x"935F" when address_in = 16#27DA# else
		x"936F" when address_in = 16#27DB# else
		x"937F" when address_in = 16#27DC# else
		x"938F" when address_in = 16#27DD# else
		x"939F" when address_in = 16#27DE# else
		x"93AF" when address_in = 16#27DF# else
		x"93BF" when address_in = 16#27E0# else
		x"93EF" when address_in = 16#27E1# else
		x"93FF" when address_in = 16#27E2# else
		x"9180" when address_in = 16#27E3# else
		x"014F" when address_in = 16#27E4# else
		x"2799" when address_in = 16#27E5# else
		x"3084" when address_in = 16#27E6# else
		x"0591" when address_in = 16#27E7# else
		x"F409" when address_in = 16#27E8# else
		x"C040" when address_in = 16#27E9# else
		x"3085" when address_in = 16#27EA# else
		x"0591" when address_in = 16#27EB# else
		x"F434" when address_in = 16#27EC# else
		x"3082" when address_in = 16#27ED# else
		x"0591" when address_in = 16#27EE# else
		x"F059" when address_in = 16#27EF# else
		x"9703" when address_in = 16#27F0# else
		x"F161" when address_in = 16#27F1# else
		x"C1D1" when address_in = 16#27F2# else
		x"3085" when address_in = 16#27F3# else
		x"0591" when address_in = 16#27F4# else
		x"F409" when address_in = 16#27F5# else
		x"C1BC" when address_in = 16#27F6# else
		x"9706" when address_in = 16#27F7# else
		x"F409" when address_in = 16#27F8# else
		x"C1C1" when address_in = 16#27F9# else
		x"C1C9" when address_in = 16#27FA# else
		x"9190" when address_in = 16#27FB# else
		x"015A" when address_in = 16#27FC# else
		x"FF97" when address_in = 16#27FD# else
		x"C002" when address_in = 16#27FE# else
		x"E081" when address_in = 16#27FF# else
		x"C001" when address_in = 16#2800# else
		x"E085" when address_in = 16#2801# else
		x"B98C" when address_in = 16#2802# else
		x"E086" when address_in = 16#2803# else
		x"9380" when address_in = 16#2804# else
		x"0151" when address_in = 16#2805# else
		x"E083" when address_in = 16#2806# else
		x"9380" when address_in = 16#2807# else
		x"014F" when address_in = 16#2808# else
		x"FF97" when address_in = 16#2809# else
		x"C1C8" when address_in = 16#280A# else
		x"E2EC" when address_in = 16#280B# else
		x"E0F9" when address_in = 16#280C# else
		x"95C8" when address_in = 16#280D# else
		x"2D80" when address_in = 16#280E# else
		x"2F28" when address_in = 16#280F# else
		x"2733" when address_in = 16#2810# else
		x"9631" when address_in = 16#2811# else
		x"95C8" when address_in = 16#2812# else
		x"2D80" when address_in = 16#2813# else
		x"2799" when address_in = 16#2814# else
		x"2F98" when address_in = 16#2815# else
		x"2788" when address_in = 16#2816# else
		x"2B28" when address_in = 16#2817# else
		x"2B39" when address_in = 16#2818# else
		x"9330" when address_in = 16#2819# else
		x"0157" when address_in = 16#281A# else
		x"9320" when address_in = 16#281B# else
		x"0156" when address_in = 16#281C# else
		x"C1B5" when address_in = 16#281D# else
		x"E084" when address_in = 16#281E# else
		x"9380" when address_in = 16#281F# else
		x"014F" when address_in = 16#2820# else
		x"9180" when address_in = 16#2821# else
		x"015A" when address_in = 16#2822# else
		x"FF87" when address_in = 16#2823# else
		x"C002" when address_in = 16#2824# else
		x"E087" when address_in = 16#2825# else
		x"C001" when address_in = 16#2826# else
		x"E082" when address_in = 16#2827# else
		x"9380" when address_in = 16#2828# else
		x"0150" when address_in = 16#2829# else
		x"9180" when address_in = 16#282A# else
		x"0150" when address_in = 16#282B# else
		x"2799" when address_in = 16#282C# else
		x"3088" when address_in = 16#282D# else
		x"0591" when address_in = 16#282E# else
		x"F409" when address_in = 16#282F# else
		x"C077" when address_in = 16#2830# else
		x"3089" when address_in = 16#2831# else
		x"0591" when address_in = 16#2832# else
		x"F43C" when address_in = 16#2833# else
		x"3082" when address_in = 16#2834# else
		x"0591" when address_in = 16#2835# else
		x"F409" when address_in = 16#2836# else
		x"C070" when address_in = 16#2837# else
		x"9707" when address_in = 16#2838# else
		x"F049" when address_in = 16#2839# else
		x"C198" when address_in = 16#283A# else
		x"3089" when address_in = 16#283B# else
		x"0591" when address_in = 16#283C# else
		x"F409" when address_in = 16#283D# else
		x"C0CF" when address_in = 16#283E# else
		x"970A" when address_in = 16#283F# else
		x"F409" when address_in = 16#2840# else
		x"C11E" when address_in = 16#2841# else
		x"C190" when address_in = 16#2842# else
		x"9170" when address_in = 16#2843# else
		x"0159" when address_in = 16#2844# else
		x"91A0" when address_in = 16#2845# else
		x"0152" when address_in = 16#2846# else
		x"91B0" when address_in = 16#2847# else
		x"0153" when address_in = 16#2848# else
		x"2FFB" when address_in = 16#2849# else
		x"2FEA" when address_in = 16#284A# else
		x"0FE7" when address_in = 16#284B# else
		x"1DF1" when address_in = 16#284C# else
		x"8160" when address_in = 16#284D# else
		x"9180" when address_in = 16#284E# else
		x"015A" when address_in = 16#284F# else
		x"FF87" when address_in = 16#2850# else
		x"C023" when address_in = 16#2851# else
		x"9180" when address_in = 16#2852# else
		x"0151" when address_in = 16#2853# else
		x"3086" when address_in = 16#2854# else
		x"F4F9" when address_in = 16#2855# else
		x"9140" when address_in = 16#2856# else
		x"0156" when address_in = 16#2857# else
		x"9150" when address_in = 16#2858# else
		x"0157" when address_in = 16#2859# else
		x"2FE5" when address_in = 16#285A# else
		x"27FF" when address_in = 16#285B# else
		x"2F86" when address_in = 16#285C# else
		x"2799" when address_in = 16#285D# else
		x"27E8" when address_in = 16#285E# else
		x"27F9" when address_in = 16#285F# else
		x"0FEE" when address_in = 16#2860# else
		x"1FFF" when address_in = 16#2861# else
		x"5DE6" when address_in = 16#2862# else
		x"4FF6" when address_in = 16#2863# else
		x"95C8" when address_in = 16#2864# else
		x"2D80" when address_in = 16#2865# else
		x"2F28" when address_in = 16#2866# else
		x"2733" when address_in = 16#2867# else
		x"9631" when address_in = 16#2868# else
		x"95C8" when address_in = 16#2869# else
		x"2D80" when address_in = 16#286A# else
		x"2784" when address_in = 16#286B# else
		x"2799" when address_in = 16#286C# else
		x"2F98" when address_in = 16#286D# else
		x"2788" when address_in = 16#286E# else
		x"2B28" when address_in = 16#286F# else
		x"2B39" when address_in = 16#2870# else
		x"9330" when address_in = 16#2871# else
		x"0157" when address_in = 16#2872# else
		x"9320" when address_in = 16#2873# else
		x"0156" when address_in = 16#2874# else
		x"9190" when address_in = 16#2875# else
		x"0151" when address_in = 16#2876# else
		x"3097" when address_in = 16#2877# else
		x"F441" when address_in = 16#2878# else
		x"E280" when address_in = 16#2879# else
		x"2768" when address_in = 16#287A# else
		x"B96C" when address_in = 16#287B# else
		x"9180" when address_in = 16#287C# else
		x"014B" when address_in = 16#287D# else
		x"9380" when address_in = 16#287E# else
		x"0151" when address_in = 16#287F# else
		x"C00F" when address_in = 16#2880# else
		x"2F86" when address_in = 16#2881# else
		x"578D" when address_in = 16#2882# else
		x"3082" when address_in = 16#2883# else
		x"F010" when address_in = 16#2884# else
		x"3063" when address_in = 16#2885# else
		x"F441" when address_in = 16#2886# else
		x"9390" when address_in = 16#2887# else
		x"014B" when address_in = 16#2888# else
		x"E087" when address_in = 16#2889# else
		x"9380" when address_in = 16#288A# else
		x"0151" when address_in = 16#288B# else
		x"E78D" when address_in = 16#288C# else
		x"B98C" when address_in = 16#288D# else
		x"C004" when address_in = 16#288E# else
		x"B96C" when address_in = 16#288F# else
		x"5F7F" when address_in = 16#2890# else
		x"9370" when address_in = 16#2891# else
		x"0159" when address_in = 16#2892# else
		x"9190" when address_in = 16#2893# else
		x"0159" when address_in = 16#2894# else
		x"3098" when address_in = 16#2895# else
		x"F009" when address_in = 16#2896# else
		x"C13B" when address_in = 16#2897# else
		x"9180" when address_in = 16#2898# else
		x"0151" when address_in = 16#2899# else
		x"3087" when address_in = 16#289A# else
		x"F409" when address_in = 16#289B# else
		x"C136" when address_in = 16#289C# else
		x"9210" when address_in = 16#289D# else
		x"0159" when address_in = 16#289E# else
		x"2FFB" when address_in = 16#289F# else
		x"2FEA" when address_in = 16#28A0# else
		x"8187" when address_in = 16#28A1# else
		x"2388" when address_in = 16#28A2# else
		x"F409" when address_in = 16#28A3# else
		x"C05F" when address_in = 16#28A4# else
		x"9390" when address_in = 16#28A5# else
		x"0150" when address_in = 16#28A6# else
		x"C12B" when address_in = 16#28A7# else
		x"9170" when address_in = 16#28A8# else
		x"0159" when address_in = 16#28A9# else
		x"91E0" when address_in = 16#28AA# else
		x"0154" when address_in = 16#28AB# else
		x"91F0" when address_in = 16#28AC# else
		x"0155" when address_in = 16#28AD# else
		x"0FE7" when address_in = 16#28AE# else
		x"1DF1" when address_in = 16#28AF# else
		x"8160" when address_in = 16#28B0# else
		x"91A0" when address_in = 16#28B1# else
		x"015A" when address_in = 16#28B2# else
		x"FFA7" when address_in = 16#28B3# else
		x"C023" when address_in = 16#28B4# else
		x"9180" when address_in = 16#28B5# else
		x"0151" when address_in = 16#28B6# else
		x"3086" when address_in = 16#28B7# else
		x"F4F9" when address_in = 16#28B8# else
		x"9140" when address_in = 16#28B9# else
		x"0156" when address_in = 16#28BA# else
		x"9150" when address_in = 16#28BB# else
		x"0157" when address_in = 16#28BC# else
		x"2FE5" when address_in = 16#28BD# else
		x"27FF" when address_in = 16#28BE# else
		x"2F86" when address_in = 16#28BF# else
		x"2799" when address_in = 16#28C0# else
		x"27E8" when address_in = 16#28C1# else
		x"27F9" when address_in = 16#28C2# else
		x"0FEE" when address_in = 16#28C3# else
		x"1FFF" when address_in = 16#28C4# else
		x"5DE6" when address_in = 16#28C5# else
		x"4FF6" when address_in = 16#28C6# else
		x"95C8" when address_in = 16#28C7# else
		x"2D80" when address_in = 16#28C8# else
		x"2F28" when address_in = 16#28C9# else
		x"2733" when address_in = 16#28CA# else
		x"9631" when address_in = 16#28CB# else
		x"95C8" when address_in = 16#28CC# else
		x"2D80" when address_in = 16#28CD# else
		x"2784" when address_in = 16#28CE# else
		x"2799" when address_in = 16#28CF# else
		x"2F98" when address_in = 16#28D0# else
		x"2788" when address_in = 16#28D1# else
		x"2B28" when address_in = 16#28D2# else
		x"2B39" when address_in = 16#28D3# else
		x"9330" when address_in = 16#28D4# else
		x"0157" when address_in = 16#28D5# else
		x"9320" when address_in = 16#28D6# else
		x"0156" when address_in = 16#28D7# else
		x"9190" when address_in = 16#28D8# else
		x"0151" when address_in = 16#28D9# else
		x"3097" when address_in = 16#28DA# else
		x"F441" when address_in = 16#28DB# else
		x"E280" when address_in = 16#28DC# else
		x"2768" when address_in = 16#28DD# else
		x"B96C" when address_in = 16#28DE# else
		x"9180" when address_in = 16#28DF# else
		x"014B" when address_in = 16#28E0# else
		x"9380" when address_in = 16#28E1# else
		x"0151" when address_in = 16#28E2# else
		x"C00F" when address_in = 16#28E3# else
		x"2F86" when address_in = 16#28E4# else
		x"578D" when address_in = 16#28E5# else
		x"3082" when address_in = 16#28E6# else
		x"F010" when address_in = 16#28E7# else
		x"3063" when address_in = 16#28E8# else
		x"F441" when address_in = 16#28E9# else
		x"9390" when address_in = 16#28EA# else
		x"014B" when address_in = 16#28EB# else
		x"E087" when address_in = 16#28EC# else
		x"9380" when address_in = 16#28ED# else
		x"0151" when address_in = 16#28EE# else
		x"E78D" when address_in = 16#28EF# else
		x"B98C" when address_in = 16#28F0# else
		x"C004" when address_in = 16#28F1# else
		x"B96C" when address_in = 16#28F2# else
		x"5F7F" when address_in = 16#28F3# else
		x"9370" when address_in = 16#28F4# else
		x"0159" when address_in = 16#28F5# else
		x"9190" when address_in = 16#28F6# else
		x"0159" when address_in = 16#28F7# else
		x"9180" when address_in = 16#28F8# else
		x"0158" when address_in = 16#28F9# else
		x"1798" when address_in = 16#28FA# else
		x"F009" when address_in = 16#28FB# else
		x"C0D6" when address_in = 16#28FC# else
		x"9180" when address_in = 16#28FD# else
		x"0151" when address_in = 16#28FE# else
		x"3087" when address_in = 16#28FF# else
		x"F409" when address_in = 16#2900# else
		x"C0D1" when address_in = 16#2901# else
		x"FFA7" when address_in = 16#2902# else
		x"C004" when address_in = 16#2903# else
		x"E089" when address_in = 16#2904# else
		x"9380" when address_in = 16#2905# else
		x"0151" when address_in = 16#2906# else
		x"C055" when address_in = 16#2907# else
		x"E086" when address_in = 16#2908# else
		x"9380" when address_in = 16#2909# else
		x"014F" when address_in = 16#290A# else
		x"E78E" when address_in = 16#290B# else
		x"B98C" when address_in = 16#290C# else
		x"C0C5" when address_in = 16#290D# else
		x"9160" when address_in = 16#290E# else
		x"0156" when address_in = 16#290F# else
		x"9180" when address_in = 16#2910# else
		x"015A" when address_in = 16#2911# else
		x"FF87" when address_in = 16#2912# else
		x"C023" when address_in = 16#2913# else
		x"9180" when address_in = 16#2914# else
		x"0151" when address_in = 16#2915# else
		x"3086" when address_in = 16#2916# else
		x"F4F9" when address_in = 16#2917# else
		x"9140" when address_in = 16#2918# else
		x"0156" when address_in = 16#2919# else
		x"9150" when address_in = 16#291A# else
		x"0157" when address_in = 16#291B# else
		x"2FE5" when address_in = 16#291C# else
		x"27FF" when address_in = 16#291D# else
		x"2F86" when address_in = 16#291E# else
		x"2799" when address_in = 16#291F# else
		x"27E8" when address_in = 16#2920# else
		x"27F9" when address_in = 16#2921# else
		x"0FEE" when address_in = 16#2922# else
		x"1FFF" when address_in = 16#2923# else
		x"5DE6" when address_in = 16#2924# else
		x"4FF6" when address_in = 16#2925# else
		x"95C8" when address_in = 16#2926# else
		x"2D80" when address_in = 16#2927# else
		x"2F28" when address_in = 16#2928# else
		x"2733" when address_in = 16#2929# else
		x"9631" when address_in = 16#292A# else
		x"95C8" when address_in = 16#292B# else
		x"2D80" when address_in = 16#292C# else
		x"2784" when address_in = 16#292D# else
		x"2799" when address_in = 16#292E# else
		x"2F98" when address_in = 16#292F# else
		x"2788" when address_in = 16#2930# else
		x"2B28" when address_in = 16#2931# else
		x"2B39" when address_in = 16#2932# else
		x"9330" when address_in = 16#2933# else
		x"0157" when address_in = 16#2934# else
		x"9320" when address_in = 16#2935# else
		x"0156" when address_in = 16#2936# else
		x"9190" when address_in = 16#2937# else
		x"0151" when address_in = 16#2938# else
		x"3097" when address_in = 16#2939# else
		x"F441" when address_in = 16#293A# else
		x"E280" when address_in = 16#293B# else
		x"2768" when address_in = 16#293C# else
		x"B96C" when address_in = 16#293D# else
		x"9180" when address_in = 16#293E# else
		x"014B" when address_in = 16#293F# else
		x"9380" when address_in = 16#2940# else
		x"0151" when address_in = 16#2941# else
		x"C00F" when address_in = 16#2942# else
		x"2F86" when address_in = 16#2943# else
		x"578D" when address_in = 16#2944# else
		x"3082" when address_in = 16#2945# else
		x"F010" when address_in = 16#2946# else
		x"3063" when address_in = 16#2947# else
		x"F441" when address_in = 16#2948# else
		x"9390" when address_in = 16#2949# else
		x"014B" when address_in = 16#294A# else
		x"E087" when address_in = 16#294B# else
		x"9380" when address_in = 16#294C# else
		x"0151" when address_in = 16#294D# else
		x"E78D" when address_in = 16#294E# else
		x"B98C" when address_in = 16#294F# else
		x"C006" when address_in = 16#2950# else
		x"B96C" when address_in = 16#2951# else
		x"9180" when address_in = 16#2952# else
		x"0159" when address_in = 16#2953# else
		x"5F8F" when address_in = 16#2954# else
		x"9380" when address_in = 16#2955# else
		x"0159" when address_in = 16#2956# else
		x"9180" when address_in = 16#2957# else
		x"0151" when address_in = 16#2958# else
		x"3087" when address_in = 16#2959# else
		x"F409" when address_in = 16#295A# else
		x"C077" when address_in = 16#295B# else
		x"E08A" when address_in = 16#295C# else
		x"9380" when address_in = 16#295D# else
		x"0150" when address_in = 16#295E# else
		x"C073" when address_in = 16#295F# else
		x"9160" when address_in = 16#2960# else
		x"0156" when address_in = 16#2961# else
		x"9170" when address_in = 16#2962# else
		x"0157" when address_in = 16#2963# else
		x"2F27" when address_in = 16#2964# else
		x"2733" when address_in = 16#2965# else
		x"2F42" when address_in = 16#2966# else
		x"9180" when address_in = 16#2967# else
		x"015A" when address_in = 16#2968# else
		x"FF87" when address_in = 16#2969# else
		x"C01D" when address_in = 16#296A# else
		x"9180" when address_in = 16#296B# else
		x"0151" when address_in = 16#296C# else
		x"3086" when address_in = 16#296D# else
		x"F4C9" when address_in = 16#296E# else
		x"2FE2" when address_in = 16#296F# else
		x"27FF" when address_in = 16#2970# else
		x"27E2" when address_in = 16#2971# else
		x"27F3" when address_in = 16#2972# else
		x"0FEE" when address_in = 16#2973# else
		x"1FFF" when address_in = 16#2974# else
		x"5DE6" when address_in = 16#2975# else
		x"4FF6" when address_in = 16#2976# else
		x"95C8" when address_in = 16#2977# else
		x"2D80" when address_in = 16#2978# else
		x"2F28" when address_in = 16#2979# else
		x"2733" when address_in = 16#297A# else
		x"9631" when address_in = 16#297B# else
		x"95C8" when address_in = 16#297C# else
		x"2D80" when address_in = 16#297D# else
		x"2786" when address_in = 16#297E# else
		x"2799" when address_in = 16#297F# else
		x"2F98" when address_in = 16#2980# else
		x"2788" when address_in = 16#2981# else
		x"2B28" when address_in = 16#2982# else
		x"2B39" when address_in = 16#2983# else
		x"9330" when address_in = 16#2984# else
		x"0157" when address_in = 16#2985# else
		x"9320" when address_in = 16#2986# else
		x"0156" when address_in = 16#2987# else
		x"9190" when address_in = 16#2988# else
		x"0151" when address_in = 16#2989# else
		x"3097" when address_in = 16#298A# else
		x"F441" when address_in = 16#298B# else
		x"E280" when address_in = 16#298C# else
		x"2748" when address_in = 16#298D# else
		x"B94C" when address_in = 16#298E# else
		x"9180" when address_in = 16#298F# else
		x"014B" when address_in = 16#2990# else
		x"9380" when address_in = 16#2991# else
		x"0151" when address_in = 16#2992# else
		x"C00F" when address_in = 16#2993# else
		x"2F84" when address_in = 16#2994# else
		x"578D" when address_in = 16#2995# else
		x"3082" when address_in = 16#2996# else
		x"F010" when address_in = 16#2997# else
		x"3043" when address_in = 16#2998# else
		x"F441" when address_in = 16#2999# else
		x"9390" when address_in = 16#299A# else
		x"014B" when address_in = 16#299B# else
		x"E087" when address_in = 16#299C# else
		x"9380" when address_in = 16#299D# else
		x"0151" when address_in = 16#299E# else
		x"E78D" when address_in = 16#299F# else
		x"B98C" when address_in = 16#29A0# else
		x"C006" when address_in = 16#29A1# else
		x"B94C" when address_in = 16#29A2# else
		x"9180" when address_in = 16#29A3# else
		x"0159" when address_in = 16#29A4# else
		x"5F8F" when address_in = 16#29A5# else
		x"9380" when address_in = 16#29A6# else
		x"0159" when address_in = 16#29A7# else
		x"9180" when address_in = 16#29A8# else
		x"0151" when address_in = 16#29A9# else
		x"3087" when address_in = 16#29AA# else
		x"F139" when address_in = 16#29AB# else
		x"E08B" when address_in = 16#29AC# else
		x"9380" when address_in = 16#29AD# else
		x"0150" when address_in = 16#29AE# else
		x"E085" when address_in = 16#29AF# else
		x"9380" when address_in = 16#29B0# else
		x"014F" when address_in = 16#29B1# else
		x"C020" when address_in = 16#29B2# else
		x"E78E" when address_in = 16#29B3# else
		x"B98C" when address_in = 16#29B4# else
		x"E086" when address_in = 16#29B5# else
		x"9380" when address_in = 16#29B6# else
		x"014F" when address_in = 16#29B7# else
		x"9210" when address_in = 16#29B8# else
		x"0150" when address_in = 16#29B9# else
		x"C018" when address_in = 16#29BA# else
		x"9856" when address_in = 16#29BB# else
		x"E081" when address_in = 16#29BC# else
		x"9380" when address_in = 16#29BD# else
		x"014F" when address_in = 16#29BE# else
		x"9210" when address_in = 16#29BF# else
		x"0151" when address_in = 16#29C0# else
		x"9180" when address_in = 16#29C1# else
		x"015A" when address_in = 16#29C2# else
		x"C00C" when address_in = 16#29C3# else
		x"9856" when address_in = 16#29C4# else
		x"9190" when address_in = 16#29C5# else
		x"015A" when address_in = 16#29C6# else
		x"6091" when address_in = 16#29C7# else
		x"9390" when address_in = 16#29C8# else
		x"015A" when address_in = 16#29C9# else
		x"E081" when address_in = 16#29CA# else
		x"9380" when address_in = 16#29CB# else
		x"014F" when address_in = 16#29CC# else
		x"9210" when address_in = 16#29CD# else
		x"0151" when address_in = 16#29CE# else
		x"2F89" when address_in = 16#29CF# else
		x"7F8E" when address_in = 16#29D0# else
		x"940E" when address_in = 16#29D1# else
		x"2D1D" when address_in = 16#29D2# else
		x"91FF" when address_in = 16#29D3# else
		x"91EF" when address_in = 16#29D4# else
		x"91BF" when address_in = 16#29D5# else
		x"91AF" when address_in = 16#29D6# else
		x"919F" when address_in = 16#29D7# else
		x"918F" when address_in = 16#29D8# else
		x"917F" when address_in = 16#29D9# else
		x"916F" when address_in = 16#29DA# else
		x"915F" when address_in = 16#29DB# else
		x"914F" when address_in = 16#29DC# else
		x"913F" when address_in = 16#29DD# else
		x"912F" when address_in = 16#29DE# else
		x"900F" when address_in = 16#29DF# else
		x"BE0F" when address_in = 16#29E0# else
		x"900F" when address_in = 16#29E1# else
		x"901F" when address_in = 16#29E2# else
		x"9518" when address_in = 16#29E3# else
		x"921F" when address_in = 16#29E4# else
		x"920F" when address_in = 16#29E5# else
		x"B60F" when address_in = 16#29E6# else
		x"920F" when address_in = 16#29E7# else
		x"2411" when address_in = 16#29E8# else
		x"92FF" when address_in = 16#29E9# else
		x"930F" when address_in = 16#29EA# else
		x"931F" when address_in = 16#29EB# else
		x"932F" when address_in = 16#29EC# else
		x"933F" when address_in = 16#29ED# else
		x"934F" when address_in = 16#29EE# else
		x"935F" when address_in = 16#29EF# else
		x"936F" when address_in = 16#29F0# else
		x"937F" when address_in = 16#29F1# else
		x"938F" when address_in = 16#29F2# else
		x"939F" when address_in = 16#29F3# else
		x"93AF" when address_in = 16#29F4# else
		x"93BF" when address_in = 16#29F5# else
		x"93CF" when address_in = 16#29F6# else
		x"93DF" when address_in = 16#29F7# else
		x"93EF" when address_in = 16#29F8# else
		x"93FF" when address_in = 16#29F9# else
		x"B0FB" when address_in = 16#29FA# else
		x"E188" when address_in = 16#29FB# else
		x"22F8" when address_in = 16#29FC# else
		x"B19C" when address_in = 16#29FD# else
		x"9180" when address_in = 16#29FE# else
		x"015B" when address_in = 16#29FF# else
		x"2F08" when address_in = 16#2A00# else
		x"2711" when address_in = 16#2A01# else
		x"3004" when address_in = 16#2A02# else
		x"0511" when address_in = 16#2A03# else
		x"F43C" when address_in = 16#2A04# else
		x"3002" when address_in = 16#2A05# else
		x"0511" when address_in = 16#2A06# else
		x"F4A4" when address_in = 16#2A07# else
		x"3001" when address_in = 16#2A08# else
		x"0511" when address_in = 16#2A09# else
		x"F051" when address_in = 16#2A0A# else
		x"C211" when address_in = 16#2A0B# else
		x"3004" when address_in = 16#2A0C# else
		x"0511" when address_in = 16#2A0D# else
		x"F409" when address_in = 16#2A0E# else
		x"C0C1" when address_in = 16#2A0F# else
		x"3005" when address_in = 16#2A10# else
		x"0511" when address_in = 16#2A11# else
		x"F409" when address_in = 16#2A12# else
		x"C1DF" when address_in = 16#2A13# else
		x"C208" when address_in = 16#2A14# else
		x"20FF" when address_in = 16#2A15# else
		x"F009" when address_in = 16#2A16# else
		x"C218" when address_in = 16#2A17# else
		x"379E" when address_in = 16#2A18# else
		x"F009" when address_in = 16#2A19# else
		x"C215" when address_in = 16#2A1A# else
		x"C013" when address_in = 16#2A1B# else
		x"20FF" when address_in = 16#2A1C# else
		x"F009" when address_in = 16#2A1D# else
		x"C1FE" when address_in = 16#2A1E# else
		x"2F89" when address_in = 16#2A1F# else
		x"2799" when address_in = 16#2A20# else
		x"3085" when address_in = 16#2A21# else
		x"0591" when address_in = 16#2A22# else
		x"F409" when address_in = 16#2A23# else
		x"C060" when address_in = 16#2A24# else
		x"3086" when address_in = 16#2A25# else
		x"0591" when address_in = 16#2A26# else
		x"F41C" when address_in = 16#2A27# else
		x"9701" when address_in = 16#2A28# else
		x"F039" when address_in = 16#2A29# else
		x"C1F2" when address_in = 16#2A2A# else
		x"378E" when address_in = 16#2A2B# else
		x"0591" when address_in = 16#2A2C# else
		x"F009" when address_in = 16#2A2D# else
		x"C1EE" when address_in = 16#2A2E# else
		x"E082" when address_in = 16#2A2F# else
		x"C1BF" when address_in = 16#2A30# else
		x"91E0" when address_in = 16#2A31# else
		x"015E" when address_in = 16#2A32# else
		x"91F0" when address_in = 16#2A33# else
		x"015F" when address_in = 16#2A34# else
		x"9730" when address_in = 16#2A35# else
		x"F439" when address_in = 16#2A36# else
		x"940E" when address_in = 16#2A37# else
		x"12DE" when address_in = 16#2A38# else
		x"9390" when address_in = 16#2A39# else
		x"015F" when address_in = 16#2A3A# else
		x"9380" when address_in = 16#2A3B# else
		x"015E" when address_in = 16#2A3C# else
		x"C01F" when address_in = 16#2A3D# else
		x"8520" when address_in = 16#2A3E# else
		x"8531" when address_in = 16#2A3F# else
		x"1521" when address_in = 16#2A40# else
		x"0531" when address_in = 16#2A41# else
		x"F0D1" when address_in = 16#2A42# else
		x"8582" when address_in = 16#2A43# else
		x"8593" when address_in = 16#2A44# else
		x"FF82" when address_in = 16#2A45# else
		x"C016" when address_in = 16#2A46# else
		x"B184" when address_in = 16#2A47# else
		x"2799" when address_in = 16#2A48# else
		x"718E" when address_in = 16#2A49# else
		x"7090" when address_in = 16#2A4A# else
		x"9595" when address_in = 16#2A4B# else
		x"9587" when address_in = 16#2A4C# else
		x"9595" when address_in = 16#2A4D# else
		x"9587" when address_in = 16#2A4E# else
		x"2F68" when address_in = 16#2A4F# else
		x"2F93" when address_in = 16#2A50# else
		x"2F82" when address_in = 16#2A51# else
		x"940E" when address_in = 16#2A52# else
		x"07EC" when address_in = 16#2A53# else
		x"91E0" when address_in = 16#2A54# else
		x"015E" when address_in = 16#2A55# else
		x"91F0" when address_in = 16#2A56# else
		x"015F" when address_in = 16#2A57# else
		x"8582" when address_in = 16#2A58# else
		x"8593" when address_in = 16#2A59# else
		x"7F8B" when address_in = 16#2A5A# else
		x"8793" when address_in = 16#2A5B# else
		x"8782" when address_in = 16#2A5C# else
		x"9180" when address_in = 16#2A5D# else
		x"015E" when address_in = 16#2A5E# else
		x"9190" when address_in = 16#2A5F# else
		x"015F" when address_in = 16#2A60# else
		x"2B89" when address_in = 16#2A61# else
		x"F409" when address_in = 16#2A62# else
		x"C1C5" when address_in = 16#2A63# else
		x"E08D" when address_in = 16#2A64# else
		x"9380" when address_in = 16#2A65# else
		x"015C" when address_in = 16#2A66# else
		x"E2EC" when address_in = 16#2A67# else
		x"E0F9" when address_in = 16#2A68# else
		x"95C8" when address_in = 16#2A69# else
		x"2D80" when address_in = 16#2A6A# else
		x"2F28" when address_in = 16#2A6B# else
		x"2733" when address_in = 16#2A6C# else
		x"9631" when address_in = 16#2A6D# else
		x"95C8" when address_in = 16#2A6E# else
		x"2D80" when address_in = 16#2A6F# else
		x"2799" when address_in = 16#2A70# else
		x"2F98" when address_in = 16#2A71# else
		x"2788" when address_in = 16#2A72# else
		x"2B28" when address_in = 16#2A73# else
		x"2B39" when address_in = 16#2A74# else
		x"9330" when address_in = 16#2A75# else
		x"0163" when address_in = 16#2A76# else
		x"9320" when address_in = 16#2A77# else
		x"0162" when address_in = 16#2A78# else
		x"9180" when address_in = 16#2A79# else
		x"0166" when address_in = 16#2A7A# else
		x"6880" when address_in = 16#2A7B# else
		x"9380" when address_in = 16#2A7C# else
		x"0166" when address_in = 16#2A7D# else
		x"9210" when address_in = 16#2A7E# else
		x"0165" when address_in = 16#2A7F# else
		x"E084" when address_in = 16#2A80# else
		x"9380" when address_in = 16#2A81# else
		x"015B" when address_in = 16#2A82# else
		x"E086" when address_in = 16#2A83# else
		x"C056" when address_in = 16#2A84# else
		x"B184" when address_in = 16#2A85# else
		x"2799" when address_in = 16#2A86# else
		x"718E" when address_in = 16#2A87# else
		x"7090" when address_in = 16#2A88# else
		x"9595" when address_in = 16#2A89# else
		x"9587" when address_in = 16#2A8A# else
		x"9595" when address_in = 16#2A8B# else
		x"9587" when address_in = 16#2A8C# else
		x"2F48" when address_in = 16#2A8D# else
		x"E462" when address_in = 16#2A8E# else
		x"E880" when address_in = 16#2A8F# else
		x"E090" when address_in = 16#2A90# else
		x"940E" when address_in = 16#2A91# else
		x"0889" when address_in = 16#2A92# else
		x"2FD9" when address_in = 16#2A93# else
		x"2FC8" when address_in = 16#2A94# else
		x"9390" when address_in = 16#2A95# else
		x"0161" when address_in = 16#2A96# else
		x"9380" when address_in = 16#2A97# else
		x"0160" when address_in = 16#2A98# else
		x"2B89" when address_in = 16#2A99# else
		x"F101" when address_in = 16#2A9A# else
		x"E083" when address_in = 16#2A9B# else
		x"9380" when address_in = 16#2A9C# else
		x"015C" when address_in = 16#2A9D# else
		x"9180" when address_in = 16#2A9E# else
		x"0166" when address_in = 16#2A9F# else
		x"FF87" when address_in = 16#2AA0# else
		x"C012" when address_in = 16#2AA1# else
		x"E3E4" when address_in = 16#2AA2# else
		x"E0F9" when address_in = 16#2AA3# else
		x"95C8" when address_in = 16#2AA4# else
		x"2D80" when address_in = 16#2AA5# else
		x"2F28" when address_in = 16#2AA6# else
		x"2733" when address_in = 16#2AA7# else
		x"9631" when address_in = 16#2AA8# else
		x"95C8" when address_in = 16#2AA9# else
		x"2D80" when address_in = 16#2AAA# else
		x"2799" when address_in = 16#2AAB# else
		x"2F98" when address_in = 16#2AAC# else
		x"2788" when address_in = 16#2AAD# else
		x"2B28" when address_in = 16#2AAE# else
		x"2B39" when address_in = 16#2AAF# else
		x"9330" when address_in = 16#2AB0# else
		x"0163" when address_in = 16#2AB1# else
		x"9320" when address_in = 16#2AB2# else
		x"0162" when address_in = 16#2AB3# else
		x"E084" when address_in = 16#2AB4# else
		x"9380" when address_in = 16#2AB5# else
		x"015B" when address_in = 16#2AB6# else
		x"E086" when address_in = 16#2AB7# else
		x"9380" when address_in = 16#2AB8# else
		x"015D" when address_in = 16#2AB9# else
		x"C013" when address_in = 16#2ABA# else
		x"9180" when address_in = 16#2ABB# else
		x"015E" when address_in = 16#2ABC# else
		x"9190" when address_in = 16#2ABD# else
		x"015F" when address_in = 16#2ABE# else
		x"9700" when address_in = 16#2ABF# else
		x"F031" when address_in = 16#2AC0# else
		x"940E" when address_in = 16#2AC1# else
		x"134D" when address_in = 16#2AC2# else
		x"93D0" when address_in = 16#2AC3# else
		x"015F" when address_in = 16#2AC4# else
		x"93C0" when address_in = 16#2AC5# else
		x"015E" when address_in = 16#2AC6# else
		x"E081" when address_in = 16#2AC7# else
		x"9380" when address_in = 16#2AC8# else
		x"015B" when address_in = 16#2AC9# else
		x"92F0" when address_in = 16#2ACA# else
		x"015C" when address_in = 16#2ACB# else
		x"92F0" when address_in = 16#2ACC# else
		x"015D" when address_in = 16#2ACD# else
		x"9210" when address_in = 16#2ACE# else
		x"0165" when address_in = 16#2ACF# else
		x"C15F" when address_in = 16#2AD0# else
		x"20FF" when address_in = 16#2AD1# else
		x"F009" when address_in = 16#2AD2# else
		x"C149" when address_in = 16#2AD3# else
		x"379D" when address_in = 16#2AD4# else
		x"F441" when address_in = 16#2AD5# else
		x"9180" when address_in = 16#2AD6# else
		x"015D" when address_in = 16#2AD7# else
		x"9380" when address_in = 16#2AD8# else
		x"014E" when address_in = 16#2AD9# else
		x"E087" when address_in = 16#2ADA# else
		x"9380" when address_in = 16#2ADB# else
		x"015D" when address_in = 16#2ADC# else
		x"C152" when address_in = 16#2ADD# else
		x"379E" when address_in = 16#2ADE# else
		x"F441" when address_in = 16#2ADF# else
		x"9180" when address_in = 16#2AE0# else
		x"015E" when address_in = 16#2AE1# else
		x"9190" when address_in = 16#2AE2# else
		x"015F" when address_in = 16#2AE3# else
		x"9700" when address_in = 16#2AE4# else
		x"F409" when address_in = 16#2AE5# else
		x"C0A5" when address_in = 16#2AE6# else
		x"C09E" when address_in = 16#2AE7# else
		x"9180" when address_in = 16#2AE8# else
		x"015D" when address_in = 16#2AE9# else
		x"3087" when address_in = 16#2AEA# else
		x"F431" when address_in = 16#2AEB# else
		x"E280" when address_in = 16#2AEC# else
		x"2798" when address_in = 16#2AED# else
		x"9180" when address_in = 16#2AEE# else
		x"014E" when address_in = 16#2AEF# else
		x"9380" when address_in = 16#2AF0# else
		x"015D" when address_in = 16#2AF1# else
		x"9180" when address_in = 16#2AF2# else
		x"015C" when address_in = 16#2AF3# else
		x"2F28" when address_in = 16#2AF4# else
		x"2733" when address_in = 16#2AF5# else
		x"302E" when address_in = 16#2AF6# else
		x"0531" when address_in = 16#2AF7# else
		x"F409" when address_in = 16#2AF8# else
		x"C09A" when address_in = 16#2AF9# else
		x"302F" when address_in = 16#2AFA# else
		x"0531" when address_in = 16#2AFB# else
		x"F444" when address_in = 16#2AFC# else
		x"3023" when address_in = 16#2AFD# else
		x"0531" when address_in = 16#2AFE# else
		x"F409" when address_in = 16#2AFF# else
		x"C093" when address_in = 16#2B00# else
		x"302D" when address_in = 16#2B01# else
		x"0531" when address_in = 16#2B02# else
		x"F051" when address_in = 16#2B03# else
		x"C118" when address_in = 16#2B04# else
		x"302F" when address_in = 16#2B05# else
		x"0531" when address_in = 16#2B06# else
		x"F409" when address_in = 16#2B07# else
		x"C0C8" when address_in = 16#2B08# else
		x"3120" when address_in = 16#2B09# else
		x"0531" when address_in = 16#2B0A# else
		x"F409" when address_in = 16#2B0B# else
		x"C0CE" when address_in = 16#2B0C# else
		x"C10F" when address_in = 16#2B0D# else
		x"91E0" when address_in = 16#2B0E# else
		x"015E" when address_in = 16#2B0F# else
		x"91F0" when address_in = 16#2B10# else
		x"015F" when address_in = 16#2B11# else
		x"379E" when address_in = 16#2B12# else
		x"F409" when address_in = 16#2B13# else
		x"C06D" when address_in = 16#2B14# else
		x"9140" when address_in = 16#2B15# else
		x"0165" when address_in = 16#2B16# else
		x"0FE4" when address_in = 16#2B17# else
		x"1DF1" when address_in = 16#2B18# else
		x"8390" when address_in = 16#2B19# else
		x"5F4F" when address_in = 16#2B1A# else
		x"9340" when address_in = 16#2B1B# else
		x"0165" when address_in = 16#2B1C# else
		x"9160" when address_in = 16#2B1D# else
		x"0162" when address_in = 16#2B1E# else
		x"9170" when address_in = 16#2B1F# else
		x"0163" when address_in = 16#2B20# else
		x"2FE7" when address_in = 16#2B21# else
		x"27FF" when address_in = 16#2B22# else
		x"2F89" when address_in = 16#2B23# else
		x"2799" when address_in = 16#2B24# else
		x"27E8" when address_in = 16#2B25# else
		x"27F9" when address_in = 16#2B26# else
		x"0FEE" when address_in = 16#2B27# else
		x"1FFF" when address_in = 16#2B28# else
		x"5DE6" when address_in = 16#2B29# else
		x"4FF6" when address_in = 16#2B2A# else
		x"95C8" when address_in = 16#2B2B# else
		x"2D80" when address_in = 16#2B2C# else
		x"2F28" when address_in = 16#2B2D# else
		x"2733" when address_in = 16#2B2E# else
		x"9631" when address_in = 16#2B2F# else
		x"95C8" when address_in = 16#2B30# else
		x"2D80" when address_in = 16#2B31# else
		x"2786" when address_in = 16#2B32# else
		x"2799" when address_in = 16#2B33# else
		x"2F98" when address_in = 16#2B34# else
		x"2788" when address_in = 16#2B35# else
		x"2B28" when address_in = 16#2B36# else
		x"2B39" when address_in = 16#2B37# else
		x"9330" when address_in = 16#2B38# else
		x"0163" when address_in = 16#2B39# else
		x"9320" when address_in = 16#2B3A# else
		x"0162" when address_in = 16#2B3B# else
		x"3048" when address_in = 16#2B3C# else
		x"F009" when address_in = 16#2B3D# else
		x"C0F1" when address_in = 16#2B3E# else
		x"91E0" when address_in = 16#2B3F# else
		x"015E" when address_in = 16#2B40# else
		x"91F0" when address_in = 16#2B41# else
		x"015F" when address_in = 16#2B42# else
		x"8127" when address_in = 16#2B43# else
		x"9320" when address_in = 16#2B44# else
		x"0164" when address_in = 16#2B45# else
		x"FD27" when address_in = 16#2B46# else
		x"C03A" when address_in = 16#2B47# else
		x"2322" when address_in = 16#2B48# else
		x"F181" when address_in = 16#2B49# else
		x"B184" when address_in = 16#2B4A# else
		x"2799" when address_in = 16#2B4B# else
		x"718E" when address_in = 16#2B4C# else
		x"7090" when address_in = 16#2B4D# else
		x"9595" when address_in = 16#2B4E# else
		x"9587" when address_in = 16#2B4F# else
		x"9595" when address_in = 16#2B50# else
		x"9587" when address_in = 16#2B51# else
		x"2F48" when address_in = 16#2B52# else
		x"E462" when address_in = 16#2B53# else
		x"2F82" when address_in = 16#2B54# else
		x"2799" when address_in = 16#2B55# else
		x"940E" when address_in = 16#2B56# else
		x"0889" when address_in = 16#2B57# else
		x"2FD9" when address_in = 16#2B58# else
		x"2FC8" when address_in = 16#2B59# else
		x"9390" when address_in = 16#2B5A# else
		x"0161" when address_in = 16#2B5B# else
		x"9380" when address_in = 16#2B5C# else
		x"0160" when address_in = 16#2B5D# else
		x"91E0" when address_in = 16#2B5E# else
		x"015E" when address_in = 16#2B5F# else
		x"91F0" when address_in = 16#2B60# else
		x"015F" when address_in = 16#2B61# else
		x"9700" when address_in = 16#2B62# else
		x"F051" when address_in = 16#2B63# else
		x"8791" when address_in = 16#2B64# else
		x"8780" when address_in = 16#2B65# else
		x"8713" when address_in = 16#2B66# else
		x"8702" when address_in = 16#2B67# else
		x"E08E" when address_in = 16#2B68# else
		x"9380" when address_in = 16#2B69# else
		x"015C" when address_in = 16#2B6A# else
		x"92F0" when address_in = 16#2B6B# else
		x"0165" when address_in = 16#2B6C# else
		x"C0C2" when address_in = 16#2B6D# else
		x"9730" when address_in = 16#2B6E# else
		x"F409" when address_in = 16#2B6F# else
		x"C0B8" when address_in = 16#2B70# else
		x"2F8E" when address_in = 16#2B71# else
		x"2F9F" when address_in = 16#2B72# else
		x"940E" when address_in = 16#2B73# else
		x"134D" when address_in = 16#2B74# else
		x"93D0" when address_in = 16#2B75# else
		x"015F" when address_in = 16#2B76# else
		x"93C0" when address_in = 16#2B77# else
		x"015E" when address_in = 16#2B78# else
		x"C0AF" when address_in = 16#2B79# else
		x"8582" when address_in = 16#2B7A# else
		x"8593" when address_in = 16#2B7B# else
		x"7F8B" when address_in = 16#2B7C# else
		x"8793" when address_in = 16#2B7D# else
		x"8782" when address_in = 16#2B7E# else
		x"8611" when address_in = 16#2B7F# else
		x"8610" when address_in = 16#2B80# else
		x"C04D" when address_in = 16#2B81# else
		x"9730" when address_in = 16#2B82# else
		x"F041" when address_in = 16#2B83# else
		x"2F8E" when address_in = 16#2B84# else
		x"2F9F" when address_in = 16#2B85# else
		x"940E" when address_in = 16#2B86# else
		x"134D" when address_in = 16#2B87# else
		x"9210" when address_in = 16#2B88# else
		x"015F" when address_in = 16#2B89# else
		x"9210" when address_in = 16#2B8A# else
		x"015E" when address_in = 16#2B8B# else
		x"E081" when address_in = 16#2B8C# else
		x"9380" when address_in = 16#2B8D# else
		x"015B" when address_in = 16#2B8E# else
		x"92F0" when address_in = 16#2B8F# else
		x"015C" when address_in = 16#2B90# else
		x"92F0" when address_in = 16#2B91# else
		x"015D" when address_in = 16#2B92# else
		x"C09C" when address_in = 16#2B93# else
		x"9180" when address_in = 16#2B94# else
		x"0165" when address_in = 16#2B95# else
		x"91E0" when address_in = 16#2B96# else
		x"0160" when address_in = 16#2B97# else
		x"91F0" when address_in = 16#2B98# else
		x"0161" when address_in = 16#2B99# else
		x"0FE8" when address_in = 16#2B9A# else
		x"1DF1" when address_in = 16#2B9B# else
		x"8390" when address_in = 16#2B9C# else
		x"5F8F" when address_in = 16#2B9D# else
		x"9380" when address_in = 16#2B9E# else
		x"0165" when address_in = 16#2B9F# else
		x"9160" when address_in = 16#2BA0# else
		x"0166" when address_in = 16#2BA1# else
		x"FF67" when address_in = 16#2BA2# else
		x"C01F" when address_in = 16#2BA3# else
		x"9140" when address_in = 16#2BA4# else
		x"0162" when address_in = 16#2BA5# else
		x"9150" when address_in = 16#2BA6# else
		x"0163" when address_in = 16#2BA7# else
		x"2FE5" when address_in = 16#2BA8# else
		x"27FF" when address_in = 16#2BA9# else
		x"2F89" when address_in = 16#2BAA# else
		x"2799" when address_in = 16#2BAB# else
		x"27E8" when address_in = 16#2BAC# else
		x"27F9" when address_in = 16#2BAD# else
		x"0FEE" when address_in = 16#2BAE# else
		x"1FFF" when address_in = 16#2BAF# else
		x"5DE6" when address_in = 16#2BB0# else
		x"4FF6" when address_in = 16#2BB1# else
		x"95C8" when address_in = 16#2BB2# else
		x"2D80" when address_in = 16#2BB3# else
		x"2F28" when address_in = 16#2BB4# else
		x"2733" when address_in = 16#2BB5# else
		x"9631" when address_in = 16#2BB6# else
		x"95C8" when address_in = 16#2BB7# else
		x"2D80" when address_in = 16#2BB8# else
		x"2784" when address_in = 16#2BB9# else
		x"2799" when address_in = 16#2BBA# else
		x"2F98" when address_in = 16#2BBB# else
		x"2788" when address_in = 16#2BBC# else
		x"2B28" when address_in = 16#2BBD# else
		x"2B39" when address_in = 16#2BBE# else
		x"9330" when address_in = 16#2BBF# else
		x"0163" when address_in = 16#2BC0# else
		x"9320" when address_in = 16#2BC1# else
		x"0162" when address_in = 16#2BC2# else
		x"9190" when address_in = 16#2BC3# else
		x"0165" when address_in = 16#2BC4# else
		x"9180" when address_in = 16#2BC5# else
		x"0164" when address_in = 16#2BC6# else
		x"1798" when address_in = 16#2BC7# else
		x"F009" when address_in = 16#2BC8# else
		x"C066" when address_in = 16#2BC9# else
		x"FF67" when address_in = 16#2BCA# else
		x"C051" when address_in = 16#2BCB# else
		x"E089" when address_in = 16#2BCC# else
		x"9380" when address_in = 16#2BCD# else
		x"015D" when address_in = 16#2BCE# else
		x"E08F" when address_in = 16#2BCF# else
		x"C007" when address_in = 16#2BD0# else
		x"2F89" when address_in = 16#2BD1# else
		x"2799" when address_in = 16#2BD2# else
		x"9390" when address_in = 16#2BD3# else
		x"014D" when address_in = 16#2BD4# else
		x"9380" when address_in = 16#2BD5# else
		x"014C" when address_in = 16#2BD6# else
		x"E180" when address_in = 16#2BD7# else
		x"9380" when address_in = 16#2BD8# else
		x"015C" when address_in = 16#2BD9# else
		x"C055" when address_in = 16#2BDA# else
		x"2F89" when address_in = 16#2BDB# else
		x"2799" when address_in = 16#2BDC# else
		x"2F38" when address_in = 16#2BDD# else
		x"2722" when address_in = 16#2BDE# else
		x"9180" when address_in = 16#2BDF# else
		x"014C" when address_in = 16#2BE0# else
		x"9190" when address_in = 16#2BE1# else
		x"014D" when address_in = 16#2BE2# else
		x"2B82" when address_in = 16#2BE3# else
		x"2B93" when address_in = 16#2BE4# else
		x"9390" when address_in = 16#2BE5# else
		x"014D" when address_in = 16#2BE6# else
		x"9380" when address_in = 16#2BE7# else
		x"014C" when address_in = 16#2BE8# else
		x"E088" when address_in = 16#2BE9# else
		x"9380" when address_in = 16#2BEA# else
		x"015D" when address_in = 16#2BEB# else
		x"E181" when address_in = 16#2BEC# else
		x"9380" when address_in = 16#2BED# else
		x"015C" when address_in = 16#2BEE# else
		x"E085" when address_in = 16#2BEF# else
		x"9380" when address_in = 16#2BF0# else
		x"015B" when address_in = 16#2BF1# else
		x"C03D" when address_in = 16#2BF2# else
		x"379E" when address_in = 16#2BF3# else
		x"F5D9" when address_in = 16#2BF4# else
		x"9210" when address_in = 16#2BF5# else
		x"015D" when address_in = 16#2BF6# else
		x"9120" when address_in = 16#2BF7# else
		x"014C" when address_in = 16#2BF8# else
		x"9130" when address_in = 16#2BF9# else
		x"014D" when address_in = 16#2BFA# else
		x"9180" when address_in = 16#2BFB# else
		x"0162" when address_in = 16#2BFC# else
		x"9190" when address_in = 16#2BFD# else
		x"0163" when address_in = 16#2BFE# else
		x"1728" when address_in = 16#2BFF# else
		x"0739" when address_in = 16#2C00# else
		x"F4B1" when address_in = 16#2C01# else
		x"91E0" when address_in = 16#2C02# else
		x"015E" when address_in = 16#2C03# else
		x"91F0" when address_in = 16#2C04# else
		x"015F" when address_in = 16#2C05# else
		x"8184" when address_in = 16#2C06# else
		x"8195" when address_in = 16#2C07# else
		x"940E" when address_in = 16#2C08# else
		x"26CA" when address_in = 16#2C09# else
		x"91E0" when address_in = 16#2C0A# else
		x"015E" when address_in = 16#2C0B# else
		x"91F0" when address_in = 16#2C0C# else
		x"015F" when address_in = 16#2C0D# else
		x"8582" when address_in = 16#2C0E# else
		x"8593" when address_in = 16#2C0F# else
		x"6099" when address_in = 16#2C10# else
		x"8793" when address_in = 16#2C11# else
		x"8782" when address_in = 16#2C12# else
		x"2F8E" when address_in = 16#2C13# else
		x"2F9F" when address_in = 16#2C14# else
		x"940E" when address_in = 16#2C15# else
		x"0EC0" when address_in = 16#2C16# else
		x"C00D" when address_in = 16#2C17# else
		x"9180" when address_in = 16#2C18# else
		x"015E" when address_in = 16#2C19# else
		x"9190" when address_in = 16#2C1A# else
		x"015F" when address_in = 16#2C1B# else
		x"C006" when address_in = 16#2C1C# else
		x"9180" when address_in = 16#2C1D# else
		x"015E" when address_in = 16#2C1E# else
		x"9190" when address_in = 16#2C1F# else
		x"015F" when address_in = 16#2C20# else
		x"9700" when address_in = 16#2C21# else
		x"F031" when address_in = 16#2C22# else
		x"940E" when address_in = 16#2C23# else
		x"134D" when address_in = 16#2C24# else
		x"9210" when address_in = 16#2C25# else
		x"015F" when address_in = 16#2C26# else
		x"9210" when address_in = 16#2C27# else
		x"015E" when address_in = 16#2C28# else
		x"E081" when address_in = 16#2C29# else
		x"9380" when address_in = 16#2C2A# else
		x"015B" when address_in = 16#2C2B# else
		x"9210" when address_in = 16#2C2C# else
		x"015C" when address_in = 16#2C2D# else
		x"9210" when address_in = 16#2C2E# else
		x"015D" when address_in = 16#2C2F# else
		x"91FF" when address_in = 16#2C30# else
		x"91EF" when address_in = 16#2C31# else
		x"91DF" when address_in = 16#2C32# else
		x"91CF" when address_in = 16#2C33# else
		x"91BF" when address_in = 16#2C34# else
		x"91AF" when address_in = 16#2C35# else
		x"919F" when address_in = 16#2C36# else
		x"918F" when address_in = 16#2C37# else
		x"917F" when address_in = 16#2C38# else
		x"916F" when address_in = 16#2C39# else
		x"915F" when address_in = 16#2C3A# else
		x"914F" when address_in = 16#2C3B# else
		x"913F" when address_in = 16#2C3C# else
		x"912F" when address_in = 16#2C3D# else
		x"911F" when address_in = 16#2C3E# else
		x"910F" when address_in = 16#2C3F# else
		x"90FF" when address_in = 16#2C40# else
		x"900F" when address_in = 16#2C41# else
		x"BE0F" when address_in = 16#2C42# else
		x"900F" when address_in = 16#2C43# else
		x"901F" when address_in = 16#2C44# else
		x"9518" when address_in = 16#2C45# else
		x"931F" when address_in = 16#2C46# else
		x"E010" when address_in = 16#2C47# else
		x"9310" when address_in = 16#2C48# else
		x"016B" when address_in = 16#2C49# else
		x"9310" when address_in = 16#2C4A# else
		x"016A" when address_in = 16#2C4B# else
		x"9310" when address_in = 16#2C4C# else
		x"0167" when address_in = 16#2C4D# else
		x"940E" when address_in = 16#2C4E# else
		x"271B" when address_in = 16#2C4F# else
		x"EF8F" when address_in = 16#2C50# else
		x"9380" when address_in = 16#2C51# else
		x"0168" when address_in = 16#2C52# else
		x"9310" when address_in = 16#2C53# else
		x"016C" when address_in = 16#2C54# else
		x"9380" when address_in = 16#2C55# else
		x"0169" when address_in = 16#2C56# else
		x"9310" when address_in = 16#2C57# else
		x"016D" when address_in = 16#2C58# else
		x"9210" when address_in = 16#2C59# else
		x"0170" when address_in = 16#2C5A# else
		x"9210" when address_in = 16#2C5B# else
		x"016F" when address_in = 16#2C5C# else
		x"E081" when address_in = 16#2C5D# else
		x"9380" when address_in = 16#2C5E# else
		x"0167" when address_in = 16#2C5F# else
		x"9380" when address_in = 16#2C60# else
		x"016B" when address_in = 16#2C61# else
		x"9380" when address_in = 16#2C62# else
		x"016A" when address_in = 16#2C63# else
		x"E080" when address_in = 16#2C64# else
		x"E090" when address_in = 16#2C65# else
		x"911F" when address_in = 16#2C66# else
		x"9508" when address_in = 16#2C67# else
		x"93CF" when address_in = 16#2C68# else
		x"93DF" when address_in = 16#2C69# else
		x"2F98" when address_in = 16#2C6A# else
		x"E0E1" when address_in = 16#2C6B# else
		x"FD66" when address_in = 16#2C6C# else
		x"E0E0" when address_in = 16#2C6D# else
		x"27FF" when address_in = 16#2C6E# else
		x"2FAE" when address_in = 16#2C6F# else
		x"2FBF" when address_in = 16#2C70# else
		x"59A9" when address_in = 16#2C71# else
		x"4FBE" when address_in = 16#2C72# else
		x"2FDB" when address_in = 16#2C73# else
		x"2FCA" when address_in = 16#2C74# else
		x"8189" when address_in = 16#2C75# else
		x"3F8F" when address_in = 16#2C76# else
		x"F041" when address_in = 16#2C77# else
		x"1789" when address_in = 16#2C78# else
		x"F419" when address_in = 16#2C79# else
		x"818B" when address_in = 16#2C7A# else
		x"3082" when address_in = 16#2C7B# else
		x"F019" when address_in = 16#2C7C# else
		x"EF80" when address_in = 16#2C7D# else
		x"EF9F" when address_in = 16#2C7E# else
		x"C00B" when address_in = 16#2C7F# else
		x"59E9" when address_in = 16#2C80# else
		x"4FFE" when address_in = 16#2C81# else
		x"8391" when address_in = 16#2C82# else
		x"E083" when address_in = 16#2C83# else
		x"9380" when address_in = 16#2C84# else
		x"0167" when address_in = 16#2C85# else
		x"8365" when address_in = 16#2C86# else
		x"E082" when address_in = 16#2C87# else
		x"8383" when address_in = 16#2C88# else
		x"E080" when address_in = 16#2C89# else
		x"E090" when address_in = 16#2C8A# else
		x"91DF" when address_in = 16#2C8B# else
		x"91CF" when address_in = 16#2C8C# else
		x"9508" when address_in = 16#2C8D# else
		x"2F28" when address_in = 16#2C8E# else
		x"3482" when address_in = 16#2C8F# else
		x"F101" when address_in = 16#2C90# else
		x"9190" when address_in = 16#2C91# else
		x"0168" when address_in = 16#2C92# else
		x"1798" when address_in = 16#2C93# else
		x"F039" when address_in = 16#2C94# else
		x"9180" when address_in = 16#2C95# else
		x"0169" when address_in = 16#2C96# else
		x"1782" when address_in = 16#2C97# else
		x"F019" when address_in = 16#2C98# else
		x"EF8F" when address_in = 16#2C99# else
		x"EF9F" when address_in = 16#2C9A# else
		x"9508" when address_in = 16#2C9B# else
		x"1792" when address_in = 16#2C9C# else
		x"F499" when address_in = 16#2C9D# else
		x"9180" when address_in = 16#2C9E# else
		x"016A" when address_in = 16#2C9F# else
		x"3081" when address_in = 16#2CA0# else
		x"F079" when address_in = 16#2CA1# else
		x"3082" when address_in = 16#2CA2# else
		x"F069" when address_in = 16#2CA3# else
		x"9180" when address_in = 16#2CA4# else
		x"0169" when address_in = 16#2CA5# else
		x"1782" when address_in = 16#2CA6# else
		x"F449" when address_in = 16#2CA7# else
		x"9180" when address_in = 16#2CA8# else
		x"016B" when address_in = 16#2CA9# else
		x"3081" when address_in = 16#2CAA# else
		x"F029" when address_in = 16#2CAB# else
		x"3082" when address_in = 16#2CAC# else
		x"F019" when address_in = 16#2CAD# else
		x"EF80" when address_in = 16#2CAE# else
		x"EF9F" when address_in = 16#2CAF# else
		x"9508" when address_in = 16#2CB0# else
		x"EF4F" when address_in = 16#2CB1# else
		x"E031" when address_in = 16#2CB2# else
		x"E6E7" when address_in = 16#2CB3# else
		x"E0F1" when address_in = 16#2CB4# else
		x"2F93" when address_in = 16#2CB5# else
		x"8181" when address_in = 16#2CB6# else
		x"1782" when address_in = 16#2CB7# else
		x"F439" when address_in = 16#2CB8# else
		x"8183" when address_in = 16#2CB9# else
		x"5081" when address_in = 16#2CBA# else
		x"3082" when address_in = 16#2CBB# else
		x"F418" when address_in = 16#2CBC# else
		x"8215" when address_in = 16#2CBD# else
		x"8341" when address_in = 16#2CBE# else
		x"8333" when address_in = 16#2CBF# else
		x"5091" when address_in = 16#2CC0# else
		x"9631" when address_in = 16#2CC1# else
		x"FF97" when address_in = 16#2CC2# else
		x"CFF2" when address_in = 16#2CC3# else
		x"9180" when address_in = 16#2CC4# else
		x"016A" when address_in = 16#2CC5# else
		x"3081" when address_in = 16#2CC6# else
		x"F431" when address_in = 16#2CC7# else
		x"9180" when address_in = 16#2CC8# else
		x"016B" when address_in = 16#2CC9# else
		x"3081" when address_in = 16#2CCA# else
		x"F411" when address_in = 16#2CCB# else
		x"9380" when address_in = 16#2CCC# else
		x"0167" when address_in = 16#2CCD# else
		x"E080" when address_in = 16#2CCE# else
		x"E090" when address_in = 16#2CCF# else
		x"9508" when address_in = 16#2CD0# else
		x"2FF9" when address_in = 16#2CD1# else
		x"2FE8" when address_in = 16#2CD2# else
		x"9120" when address_in = 16#2CD3# else
		x"016A" when address_in = 16#2CD4# else
		x"3021" when address_in = 16#2CD5# else
		x"F419" when address_in = 16#2CD6# else
		x"EE8A" when address_in = 16#2CD7# else
		x"EF9F" when address_in = 16#2CD8# else
		x"9508" when address_in = 16#2CD9# else
		x"9180" when address_in = 16#2CDA# else
		x"0168" when address_in = 16#2CDB# else
		x"1784" when address_in = 16#2CDC# else
		x"F411" when address_in = 16#2CDD# else
		x"3022" when address_in = 16#2CDE# else
		x"F019" when address_in = 16#2CDF# else
		x"EF80" when address_in = 16#2CE0# else
		x"EF9F" when address_in = 16#2CE1# else
		x"9508" when address_in = 16#2CE2# else
		x"93F0" when address_in = 16#2CE3# else
		x"0170" when address_in = 16#2CE4# else
		x"93E0" when address_in = 16#2CE5# else
		x"016F" when address_in = 16#2CE6# else
		x"9140" when address_in = 16#2CE7# else
		x"016C" when address_in = 16#2CE8# else
		x"2F8E" when address_in = 16#2CE9# else
		x"2F9F" when address_in = 16#2CEA# else
		x"940E" when address_in = 16#2CEB# else
		x"2740" when address_in = 16#2CEC# else
		x"2388" when address_in = 16#2CED# else
		x"F441" when address_in = 16#2CEE# else
		x"E083" when address_in = 16#2CEF# else
		x"9380" when address_in = 16#2CF0# else
		x"016A" when address_in = 16#2CF1# else
		x"9380" when address_in = 16#2CF2# else
		x"0167" when address_in = 16#2CF3# else
		x"E080" when address_in = 16#2CF4# else
		x"E090" when address_in = 16#2CF5# else
		x"9508" when address_in = 16#2CF6# else
		x"EF80" when address_in = 16#2CF7# else
		x"EF9F" when address_in = 16#2CF8# else
		x"9508" when address_in = 16#2CF9# else
		x"2F28" when address_in = 16#2CFA# else
		x"9190" when address_in = 16#2CFB# else
		x"016B" when address_in = 16#2CFC# else
		x"3091" when address_in = 16#2CFD# else
		x"F419" when address_in = 16#2CFE# else
		x"EE8A" when address_in = 16#2CFF# else
		x"EF9F" when address_in = 16#2D00# else
		x"9508" when address_in = 16#2D01# else
		x"9180" when address_in = 16#2D02# else
		x"0169" when address_in = 16#2D03# else
		x"1786" when address_in = 16#2D04# else
		x"F411" when address_in = 16#2D05# else
		x"3092" when address_in = 16#2D06# else
		x"F019" when address_in = 16#2D07# else
		x"EF80" when address_in = 16#2D08# else
		x"EF9F" when address_in = 16#2D09# else
		x"9508" when address_in = 16#2D0A# else
		x"9160" when address_in = 16#2D0B# else
		x"016D" when address_in = 16#2D0C# else
		x"2F82" when address_in = 16#2D0D# else
		x"940E" when address_in = 16#2D0E# else
		x"2771" when address_in = 16#2D0F# else
		x"2388" when address_in = 16#2D10# else
		x"F441" when address_in = 16#2D11# else
		x"E083" when address_in = 16#2D12# else
		x"9380" when address_in = 16#2D13# else
		x"016B" when address_in = 16#2D14# else
		x"9380" when address_in = 16#2D15# else
		x"0167" when address_in = 16#2D16# else
		x"E080" when address_in = 16#2D17# else
		x"E090" when address_in = 16#2D18# else
		x"9508" when address_in = 16#2D19# else
		x"EF80" when address_in = 16#2D1A# else
		x"EF9F" when address_in = 16#2D1B# else
		x"9508" when address_in = 16#2D1C# else
		x"92EF" when address_in = 16#2D1D# else
		x"92FF" when address_in = 16#2D1E# else
		x"930F" when address_in = 16#2D1F# else
		x"931F" when address_in = 16#2D20# else
		x"2F98" when address_in = 16#2D21# else
		x"9130" when address_in = 16#2D22# else
		x"0168" when address_in = 16#2D23# else
		x"3F3F" when address_in = 16#2D24# else
		x"F0F1" when address_in = 16#2D25# else
		x"9180" when address_in = 16#2D26# else
		x"016A" when address_in = 16#2D27# else
		x"3083" when address_in = 16#2D28# else
		x"F4D1" when address_in = 16#2D29# else
		x"E082" when address_in = 16#2D2A# else
		x"9380" when address_in = 16#2D2B# else
		x"016A" when address_in = 16#2D2C# else
		x"2F89" when address_in = 16#2D2D# else
		x"2799" when address_in = 16#2D2E# else
		x"2F08" when address_in = 16#2D2F# else
		x"2F19" when address_in = 16#2D30# else
		x"7001" when address_in = 16#2D31# else
		x"7010" when address_in = 16#2D32# else
		x"FF80" when address_in = 16#2D33# else
		x"C006" when address_in = 16#2D34# else
		x"E492" when address_in = 16#2D35# else
		x"2EE9" when address_in = 16#2D36# else
		x"2CF1" when address_in = 16#2D37# else
		x"E000" when address_in = 16#2D38# else
		x"E010" when address_in = 16#2D39# else
		x"C003" when address_in = 16#2D3A# else
		x"E480" when address_in = 16#2D3B# else
		x"2EE8" when address_in = 16#2D3C# else
		x"2CF1" when address_in = 16#2D3D# else
		x"E020" when address_in = 16#2D3E# else
		x"E442" when address_in = 16#2D3F# else
		x"2F64" when address_in = 16#2D40# else
		x"2F83" when address_in = 16#2D41# else
		x"940E" when address_in = 16#2D42# else
		x"0FD8" when address_in = 16#2D43# else
		x"911F" when address_in = 16#2D44# else
		x"910F" when address_in = 16#2D45# else
		x"90FF" when address_in = 16#2D46# else
		x"90EF" when address_in = 16#2D47# else
		x"9508" when address_in = 16#2D48# else
		x"92EF" when address_in = 16#2D49# else
		x"92FF" when address_in = 16#2D4A# else
		x"930F" when address_in = 16#2D4B# else
		x"931F" when address_in = 16#2D4C# else
		x"FF60" when address_in = 16#2D4D# else
		x"C00E" when address_in = 16#2D4E# else
		x"9180" when address_in = 16#2D4F# else
		x"0169" when address_in = 16#2D50# else
		x"3F8F" when address_in = 16#2D51# else
		x"F051" when address_in = 16#2D52# else
		x"E420" when address_in = 16#2D53# else
		x"2EE2" when address_in = 16#2D54# else
		x"2CF1" when address_in = 16#2D55# else
		x"E000" when address_in = 16#2D56# else
		x"E010" when address_in = 16#2D57# else
		x"E020" when address_in = 16#2D58# else
		x"E04F" when address_in = 16#2D59# else
		x"E462" when address_in = 16#2D5A# else
		x"940E" when address_in = 16#2D5B# else
		x"0FD8" when address_in = 16#2D5C# else
		x"911F" when address_in = 16#2D5D# else
		x"910F" when address_in = 16#2D5E# else
		x"90FF" when address_in = 16#2D5F# else
		x"90EF" when address_in = 16#2D60# else
		x"9508" when address_in = 16#2D61# else
		x"2F38" when address_in = 16#2D62# else
		x"2F96" when address_in = 16#2D63# else
		x"B72F" when address_in = 16#2D64# else
		x"94F8" when address_in = 16#2D65# else
		x"7097" when address_in = 16#2D66# else
		x"6098" when address_in = 16#2D67# else
		x"BE17" when address_in = 16#2D68# else
		x"B780" when address_in = 16#2D69# else
		x"6088" when address_in = 16#2D6A# else
		x"BF80" when address_in = 16#2D6B# else
		x"BF93" when address_in = 16#2D6C# else
		x"BE12" when address_in = 16#2D6D# else
		x"BF31" when address_in = 16#2D6E# else
		x"B787" when address_in = 16#2D6F# else
		x"6082" when address_in = 16#2D70# else
		x"BF87" when address_in = 16#2D71# else
		x"BF2F" when address_in = 16#2D72# else
		x"940E" when address_in = 16#2D73# else
		x"1B5A" when address_in = 16#2D74# else
		x"9508" when address_in = 16#2D75# else
		x"2F26" when address_in = 16#2D76# else
		x"2F37" when address_in = 16#2D77# else
		x"2F48" when address_in = 16#2D78# else
		x"2F59" when address_in = 16#2D79# else
		x"B780" when address_in = 16#2D7A# else
		x"2799" when address_in = 16#2D7B# else
		x"7086" when address_in = 16#2D7C# else
		x"7090" when address_in = 16#2D7D# else
		x"2B89" when address_in = 16#2D7E# else
		x"F7D1" when address_in = 16#2D7F# else
		x"3F2B" when address_in = 16#2D80# else
		x"0531" when address_in = 16#2D81# else
		x"0541" when address_in = 16#2D82# else
		x"0551" when address_in = 16#2D83# else
		x"F014" when address_in = 16#2D84# else
		x"EF6A" when address_in = 16#2D85# else
		x"C009" when address_in = 16#2D86# else
		x"3023" when address_in = 16#2D87# else
		x"0531" when address_in = 16#2D88# else
		x"0541" when address_in = 16#2D89# else
		x"0551" when address_in = 16#2D8A# else
		x"F414" when address_in = 16#2D8B# else
		x"E062" when address_in = 16#2D8C# else
		x"C002" when address_in = 16#2D8D# else
		x"2F62" when address_in = 16#2D8E# else
		x"5061" when address_in = 16#2D8F# else
		x"BE12" when address_in = 16#2D90# else
		x"BF61" when address_in = 16#2D91# else
		x"9508" when address_in = 16#2D92# else
		x"E980" when address_in = 16#2D93# else
		x"E09A" when address_in = 16#2D94# else
		x"B983" when address_in = 16#2D95# else
		x"2F89" when address_in = 16#2D96# else
		x"2799" when address_in = 16#2D97# else
		x"B982" when address_in = 16#2D98# else
		x"E880" when address_in = 16#2D99# else
		x"E090" when address_in = 16#2D9A# else
		x"BB8C" when address_in = 16#2D9B# else
		x"BA1F" when address_in = 16#2D9C# else
		x"9508" when address_in = 16#2D9D# else
		x"FD87" when address_in = 16#2D9E# else
		x"C002" when address_in = 16#2D9F# else
		x"E087" when address_in = 16#2DA0# else
		x"C019" when address_in = 16#2DA1# else
		x"940E" when address_in = 16#2DA2# else
		x"0B28" when address_in = 16#2DA3# else
		x"2FF9" when address_in = 16#2DA4# else
		x"2FE8" when address_in = 16#2DA5# else
		x"2B89" when address_in = 16#2DA6# else
		x"F419" when address_in = 16#2DA7# else
		x"EE8A" when address_in = 16#2DA8# else
		x"EF9F" when address_in = 16#2DA9# else
		x"9508" when address_in = 16#2DAA# else
		x"8182" when address_in = 16#2DAB# else
		x"8193" when address_in = 16#2DAC# else
		x"27AA" when address_in = 16#2DAD# else
		x"27BB" when address_in = 16#2DAE# else
		x"0F88" when address_in = 16#2DAF# else
		x"1F99" when address_in = 16#2DB0# else
		x"1FAA" when address_in = 16#2DB1# else
		x"1FBB" when address_in = 16#2DB2# else
		x"960A" when address_in = 16#2DB3# else
		x"1DA1" when address_in = 16#2DB4# else
		x"1DB1" when address_in = 16#2DB5# else
		x"BFAB" when address_in = 16#2DB6# else
		x"2FF9" when address_in = 16#2DB7# else
		x"2FE8" when address_in = 16#2DB8# else
		x"95D8" when address_in = 16#2DB9# else
		x"2D80" when address_in = 16#2DBA# else
		x"2799" when address_in = 16#2DBB# else
		x"FD87" when address_in = 16#2DBC# else
		x"9590" when address_in = 16#2DBD# else
		x"9508" when address_in = 16#2DBE# else
		x"931F" when address_in = 16#2DBF# else
		x"93CF" when address_in = 16#2DC0# else
		x"93DF" when address_in = 16#2DC1# else
		x"E081" when address_in = 16#2DC2# else
		x"940E" when address_in = 16#2DC3# else
		x"26CF" when address_in = 16#2DC4# else
		x"E085" when address_in = 16#2DC5# else
		x"940E" when address_in = 16#2DC6# else
		x"26CF" when address_in = 16#2DC7# else
		x"E086" when address_in = 16#2DC8# else
		x"940E" when address_in = 16#2DC9# else
		x"26CF" when address_in = 16#2DCA# else
		x"EFCF" when address_in = 16#2DCB# else
		x"EFDF" when address_in = 16#2DCC# else
		x"E010" when address_in = 16#2DCD# else
		x"95A8" when address_in = 16#2DCE# else
		x"9720" when address_in = 16#2DCF# else
		x"F511" when address_in = 16#2DD0# else
		x"2F81" when address_in = 16#2DD1# else
		x"2799" when address_in = 16#2DD2# else
		x"3081" when address_in = 16#2DD3# else
		x"0591" when address_in = 16#2DD4# else
		x"F071" when address_in = 16#2DD5# else
		x"3082" when address_in = 16#2DD6# else
		x"0591" when address_in = 16#2DD7# else
		x"F41C" when address_in = 16#2DD8# else
		x"2B89" when address_in = 16#2DD9# else
		x"F021" when address_in = 16#2DDA# else
		x"C013" when address_in = 16#2DDB# else
		x"9702" when address_in = 16#2DDC# else
		x"F059" when address_in = 16#2DDD# else
		x"C010" when address_in = 16#2DDE# else
		x"E087" when address_in = 16#2DDF# else
		x"940E" when address_in = 16#2DE0# else
		x"26CF" when address_in = 16#2DE1# else
		x"E088" when address_in = 16#2DE2# else
		x"C009" when address_in = 16#2DE3# else
		x"E088" when address_in = 16#2DE4# else
		x"940E" when address_in = 16#2DE5# else
		x"26CF" when address_in = 16#2DE6# else
		x"E089" when address_in = 16#2DE7# else
		x"C004" when address_in = 16#2DE8# else
		x"E089" when address_in = 16#2DE9# else
		x"940E" when address_in = 16#2DEA# else
		x"26CF" when address_in = 16#2DEB# else
		x"E087" when address_in = 16#2DEC# else
		x"940E" when address_in = 16#2DED# else
		x"26CF" when address_in = 16#2DEE# else
		x"5F1F" when address_in = 16#2DEF# else
		x"3013" when address_in = 16#2DF0# else
		x"F409" when address_in = 16#2DF1# else
		x"E010" when address_in = 16#2DF2# else
		x"9721" when address_in = 16#2DF3# else
		x"CFD9" when address_in = 16#2DF4# else
		x"FF80" when address_in = 16#2DF5# else
		x"C002" when address_in = 16#2DF6# else
		x"98D8" when address_in = 16#2DF7# else
		x"C001" when address_in = 16#2DF8# else
		x"9AD8" when address_in = 16#2DF9# else
		x"9586" when address_in = 16#2DFA# else
		x"FF80" when address_in = 16#2DFB# else
		x"C002" when address_in = 16#2DFC# else
		x"98D9" when address_in = 16#2DFD# else
		x"C001" when address_in = 16#2DFE# else
		x"9AD9" when address_in = 16#2DFF# else
		x"9586" when address_in = 16#2E00# else
		x"FF80" when address_in = 16#2E01# else
		x"C002" when address_in = 16#2E02# else
		x"98DA" when address_in = 16#2E03# else
		x"9508" when address_in = 16#2E04# else
		x"9ADA" when address_in = 16#2E05# else
		x"9508" when address_in = 16#2E06# else
		x"931F" when address_in = 16#2E07# else
		x"93CF" when address_in = 16#2E08# else
		x"93DF" when address_in = 16#2E09# else
		x"2F18" when address_in = 16#2E0A# else
		x"EFCF" when address_in = 16#2E0B# else
		x"EFDF" when address_in = 16#2E0C# else
		x"940E" when address_in = 16#2E0D# else
		x"2DF5" when address_in = 16#2E0E# else
		x"E080" when address_in = 16#2E0F# else
		x"95A8" when address_in = 16#2E10# else
		x"9720" when address_in = 16#2E11# else
		x"F451" when address_in = 16#2E12# else
		x"2388" when address_in = 16#2E13# else
		x"F029" when address_in = 16#2E14# else
		x"2F81" when address_in = 16#2E15# else
		x"940E" when address_in = 16#2E16# else
		x"2DF5" when address_in = 16#2E17# else
		x"E080" when address_in = 16#2E18# else
		x"C003" when address_in = 16#2E19# else
		x"940E" when address_in = 16#2E1A# else
		x"2DF5" when address_in = 16#2E1B# else
		x"E081" when address_in = 16#2E1C# else
		x"9721" when address_in = 16#2E1D# else
		x"CFF1" when address_in = 16#2E1E# else
		x"921F" when address_in = 16#2E1F# else
		x"920F" when address_in = 16#2E20# else
		x"B60F" when address_in = 16#2E21# else
		x"920F" when address_in = 16#2E22# else
		x"2411" when address_in = 16#2E23# else
		x"938F" when address_in = 16#2E24# else
		x"E383" when address_in = 16#2E25# else
		x"BB8B" when address_in = 16#2E26# else
		x"EF80" when address_in = 16#2E27# else
		x"BB81" when address_in = 16#2E28# else
		x"E282" when address_in = 16#2E29# else
		x"BB8B" when address_in = 16#2E2A# else
		x"CFFF" when address_in = 16#2E2B# else
		x"27AA" when address_in = 16#2E2C# else
		x"2FE8" when address_in = 16#2E2D# else
		x"2FF9" when address_in = 16#2E2E# else
		x"0FEE" when address_in = 16#2E2F# else
		x"1FFF" when address_in = 16#2E30# else
		x"1FAA" when address_in = 16#2E31# else
		x"BFAB" when address_in = 16#2E32# else
		x"95C8" when address_in = 16#2E33# else
		x"2DA0" when address_in = 16#2E34# else
		x"9631" when address_in = 16#2E35# else
		x"95C8" when address_in = 16#2E36# else
		x"2DB0" when address_in = 16#2E37# else
		x"93AF" when address_in = 16#2E38# else
		x"93BF" when address_in = 16#2E39# else
		x"9635" when address_in = 16#2E3A# else
		x"B60F" when address_in = 16#2E3B# else
		x"94F8" when address_in = 16#2E3C# else
		x"920F" when address_in = 16#2E3D# else
		x"9010" when address_in = 16#2E3E# else
		x"0173" when address_in = 16#2E3F# else
		x"91A0" when address_in = 16#2E40# else
		x"0174" when address_in = 16#2E41# else
		x"91B0" when address_in = 16#2E42# else
		x"0175" when address_in = 16#2E43# else
		x"921D" when address_in = 16#2E44# else
		x"93A0" when address_in = 16#2E45# else
		x"0174" when address_in = 16#2E46# else
		x"93B0" when address_in = 16#2E47# else
		x"0175" when address_in = 16#2E48# else
		x"95C8" when address_in = 16#2E49# else
		x"2DA0" when address_in = 16#2E4A# else
		x"3FAF" when address_in = 16#2E4B# else
		x"F411" when address_in = 16#2E4C# else
		x"91A0" when address_in = 16#2E4D# else
		x"0173" when address_in = 16#2E4E# else
		x"93A0" when address_in = 16#2E4F# else
		x"0173" when address_in = 16#2E50# else
		x"900F" when address_in = 16#2E51# else
		x"BE0F" when address_in = 16#2E52# else
		x"91FF" when address_in = 16#2E53# else
		x"91EF" when address_in = 16#2E54# else
		x"2411" when address_in = 16#2E55# else
		x"9509" when address_in = 16#2E56# else
		x"B60F" when address_in = 16#2E57# else
		x"94F8" when address_in = 16#2E58# else
		x"91A0" when address_in = 16#2E59# else
		x"0174" when address_in = 16#2E5A# else
		x"91B0" when address_in = 16#2E5B# else
		x"0175" when address_in = 16#2E5C# else
		x"901E" when address_in = 16#2E5D# else
		x"93A0" when address_in = 16#2E5E# else
		x"0174" when address_in = 16#2E5F# else
		x"93B0" when address_in = 16#2E60# else
		x"0175" when address_in = 16#2E61# else
		x"9210" when address_in = 16#2E62# else
		x"0173" when address_in = 16#2E63# else
		x"BE0F" when address_in = 16#2E64# else
		x"2411" when address_in = 16#2E65# else
		x"9508" when address_in = 16#2E66# else
		x"2FE6" when address_in = 16#2E67# else
		x"2FF7" when address_in = 16#2E68# else
		x"2FA8" when address_in = 16#2E69# else
		x"2FB9" when address_in = 16#2E6A# else
		x"FF40" when address_in = 16#2E6B# else
		x"C005" when address_in = 16#2E6C# else
		x"C002" when address_in = 16#2E6D# else
		x"9001" when address_in = 16#2E6E# else
		x"920D" when address_in = 16#2E6F# else
		x"9001" when address_in = 16#2E70# else
		x"920D" when address_in = 16#2E71# else
		x"5042" when address_in = 16#2E72# else
		x"4050" when address_in = 16#2E73# else
		x"F7C8" when address_in = 16#2E74# else
		x"9508" when address_in = 16#2E75# else
		x"2755" when address_in = 16#2E76# else
		x"2400" when address_in = 16#2E77# else
		x"FF80" when address_in = 16#2E78# else
		x"C002" when address_in = 16#2E79# else
		x"0E06" when address_in = 16#2E7A# else
		x"1F57" when address_in = 16#2E7B# else
		x"0F66" when address_in = 16#2E7C# else
		x"1F77" when address_in = 16#2E7D# else
		x"1561" when address_in = 16#2E7E# else
		x"0571" when address_in = 16#2E7F# else
		x"F021" when address_in = 16#2E80# else
		x"9596" when address_in = 16#2E81# else
		x"9587" when address_in = 16#2E82# else
		x"9700" when address_in = 16#2E83# else
		x"F799" when address_in = 16#2E84# else
		x"2F95" when address_in = 16#2E85# else
		x"2D80" when address_in = 16#2E86# else
		x"9508" when address_in = 16#2E87# else
		x"27FF" when address_in = 16#2E88# else
		x"27EE" when address_in = 16#2E89# else
		x"27BB" when address_in = 16#2E8A# else
		x"27AA" when address_in = 16#2E8B# else
		x"FF60" when address_in = 16#2E8C# else
		x"C004" when address_in = 16#2E8D# else
		x"0FA2" when address_in = 16#2E8E# else
		x"1FB3" when address_in = 16#2E8F# else
		x"1FE4" when address_in = 16#2E90# else
		x"1FF5" when address_in = 16#2E91# else
		x"0F22" when address_in = 16#2E92# else
		x"1F33" when address_in = 16#2E93# else
		x"1F44" when address_in = 16#2E94# else
		x"1F55" when address_in = 16#2E95# else
		x"9596" when address_in = 16#2E96# else
		x"9587" when address_in = 16#2E97# else
		x"9577" when address_in = 16#2E98# else
		x"9567" when address_in = 16#2E99# else
		x"F789" when address_in = 16#2E9A# else
		x"9700" when address_in = 16#2E9B# else
		x"0776" when address_in = 16#2E9C# else
		x"F771" when address_in = 16#2E9D# else
		x"2F9F" when address_in = 16#2E9E# else
		x"2F8E" when address_in = 16#2E9F# else
		x"2F7B" when address_in = 16#2EA0# else
		x"2F6A" when address_in = 16#2EA1# else
		x"9508" when address_in = 16#2EA2# else
		x"CFFF" when address_in = 16#2EA3# else
		x"ffff";
end rtl;
